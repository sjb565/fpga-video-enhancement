`timescale 1ns / 1ps
`default_nettype none

module kernel_4_tb;

    //make logics for inputs and outputs!
    logic clk_in;
    logic rst_in;
    logic valid_in;
    logic [5:0] pixel_array_in [3:0][3:0];
    logic [8:0] pixel_out;

    kernel_4 uut (
        .clk_in(clk_in),
        .p(pixel_array_in),
        .pixel_out(pixel_out)
    );
    always begin
        #5;  //every 5 ns switch...so period of clock is 10 ns...100 MHz clock
        clk_in = !clk_in;
    end

    //initial block...this is our test simulation
    initial begin
        
		$dumpfile("test/kernel_4.vcd"); //file to store value change dump (vcd)
		$dumpvars(0,kernel_4_tb); //store everything at the current level and below
		$display("Starting Sim"); //print nice message
		clk_in = 0; //initialize clk (super important)
		rst_in = 0; //initialize rst (super important)
		
		#10;  //wait a little bit of time at beginning
		rst_in = 1; //reset system
		#10; //hold high for a few clock cycles
		rst_in=0;
		
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 0;
		#10;
		
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 32;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 32;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 32;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 32;
		#10;
		
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 63;
		#10;
		
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 63;
		#10;
		
		$display("Input: \n[[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0]]");
		$display("Expect: 0, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Input: \n[[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32]]");
		$display("Expect: 128, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 43;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 13;
		pixel_array_in[1][2] = 1;
		pixel_array_in[1][3] = 9;
		pixel_array_in[2][0] = 20;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 36;
		pixel_array_in[2][3] = 26;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 60;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 9;
		#10;
		
		$display("Input: \n[[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63]]");
		$display("Expect: 252, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 10;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 40;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 5;
		pixel_array_in[1][2] = 14;
		pixel_array_in[1][3] = 21;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 46;
		pixel_array_in[2][2] = 39;
		pixel_array_in[2][3] = 57;
		pixel_array_in[3][0] = 9;
		pixel_array_in[3][1] = 16;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 31;
		#10;
		
		$display("Input: \n[[63, 0, 0, 63],\n[0, 63, 63, 0],\n[0, 63, 63, 0],\n[63, 0, 0, 63]]");
		$display("Expect: 384>val>255, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 62;
		pixel_array_in[0][1] = 49;
		pixel_array_in[0][2] = 3;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 26;
		pixel_array_in[1][1] = 41;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 50;
		pixel_array_in[2][0] = 3;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 34;
		pixel_array_in[2][3] = 40;
		pixel_array_in[3][0] = 3;
		pixel_array_in[3][1] = 8;
		pixel_array_in[3][2] = 40;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[0, 63, 63, 0],\n[63, 0, 0, 63],\n[63, 0, 0, 63],\n[0, 63, 63, 0]]");
		$display("Expect: val>383, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 6;
		pixel_array_in[0][1] = 43;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 26;
		pixel_array_in[2][0] = 51;
		pixel_array_in[2][1] = 62;
		pixel_array_in[2][2] = 46;
		pixel_array_in[2][3] = 47;
		pixel_array_in[3][0] = 7;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[57, 0, 52, 43],\n[10, 13, 1, 9],\n[20, 11, 36, 26],\n[61, 60, 60, 9]]");
		$display("Expect: 42, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 62;
		pixel_array_in[0][1] = 46;
		pixel_array_in[0][2] = 3;
		pixel_array_in[0][3] = 48;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 51;
		pixel_array_in[1][2] = 18;
		pixel_array_in[1][3] = 59;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 8;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 61;
		pixel_array_in[3][2] = 49;
		pixel_array_in[3][3] = 51;
		#10;
		
		$display("Input: \n[[10, 19, 40, 58],\n[13, 5, 14, 21],\n[40, 46, 39, 57],\n[9, 16, 27, 31]]");
		$display("Expect: 103, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 60;
		pixel_array_in[0][1] = 51;
		pixel_array_in[0][2] = 39;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 17;
		pixel_array_in[1][1] = 14;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 52;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 14;
		pixel_array_in[3][1] = 7;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 59;
		#10;
		
		$display("Input: \n[[62, 49, 3, 15],\n[26, 41, 15, 50],\n[3, 11, 34, 40],\n[3, 8, 40, 60]]");
		$display("Expect: 103, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 14;
		pixel_array_in[0][1] = 61;
		pixel_array_in[0][2] = 26;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 37;
		pixel_array_in[1][1] = 43;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 43;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 46;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 37;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 9;
		#10;
		
		$display("Input: \n[[6, 43, 48, 58],\n[47, 27, 22, 26],\n[51, 62, 46, 47],\n[7, 48, 48, 7]]");
		$display("Expect: 164, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 53;
		pixel_array_in[0][2] = 59;
		pixel_array_in[0][3] = 35;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 58;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 61;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 58;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[62, 46, 3, 48],\n[0, 51, 18, 59],\n[31, 32, 8, 18],\n[25, 61, 49, 51]]");
		$display("Expect: 142, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 56;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 36;
		pixel_array_in[1][1] = 29;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 19;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 61;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 12;
		pixel_array_in[3][0] = 54;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 5;
		pixel_array_in[3][3] = 51;
		#10;
		
		$display("Input: \n[[60, 51, 39, 53],\n[17, 14, 56, 56],\n[52, 0, 22, 41],\n[14, 7, 32, 59]]");
		$display("Expect: 36, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 20;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 1;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 10;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 44;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 20;
		pixel_array_in[3][3] = 25;
		#10;
		
		$display("Input: \n[[14, 61, 26, 58],\n[37, 43, 13, 43],\n[12, 46, 62, 43],\n[37, 59, 61, 9]]");
		$display("Expect: 169, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 46;
		pixel_array_in[0][1] = 42;
		pixel_array_in[0][2] = 41;
		pixel_array_in[0][3] = 49;
		pixel_array_in[1][0] = 41;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 51;
		pixel_array_in[1][3] = 55;
		pixel_array_in[2][0] = 2;
		pixel_array_in[2][1] = 48;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 52;
		pixel_array_in[3][0] = 11;
		pixel_array_in[3][1] = 41;
		pixel_array_in[3][2] = 14;
		pixel_array_in[3][3] = 37;
		#10;
		
		$display("Input: \n[[21, 53, 59, 35],\n[22, 58, 11, 0],\n[30, 36, 30, 61],\n[40, 0, 58, 2]]");
		$display("Expect: 176, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 17;
		pixel_array_in[0][1] = 16;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 14;
		pixel_array_in[1][1] = 6;
		pixel_array_in[1][2] = 27;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 14;
		pixel_array_in[2][2] = 3;
		pixel_array_in[2][3] = 26;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 32;
		#10;
		
		$display("Input: \n[[8, 17, 56, 55],\n[36, 29, 37, 19],\n[1, 61, 43, 12],\n[54, 59, 5, 51]]");
		$display("Expect: 190, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 4;
		pixel_array_in[1][0] = 42;
		pixel_array_in[1][1] = 4;
		pixel_array_in[1][2] = 35;
		pixel_array_in[1][3] = 30;
		pixel_array_in[2][0] = 23;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 24;
		pixel_array_in[2][3] = 51;
		pixel_array_in[3][0] = 7;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 5;
		#10;
		
		$display("Input: \n[[21, 25, 0, 33],\n[28, 20, 50, 1],\n[40, 1, 10, 0],\n[44, 55, 20, 25]]");
		$display("Expect: 43, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 11;
		pixel_array_in[0][1] = 13;
		pixel_array_in[0][2] = 47;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 35;
		pixel_array_in[1][1] = 15;
		pixel_array_in[1][2] = 57;
		pixel_array_in[1][3] = 8;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 27;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 40;
		pixel_array_in[3][0] = 58;
		pixel_array_in[3][1] = 43;
		pixel_array_in[3][2] = 26;
		pixel_array_in[3][3] = 43;
		#10;
		
		$display("Input: \n[[46, 42, 41, 49],\n[41, 1, 51, 55],\n[2, 48, 52, 52],\n[11, 41, 14, 37]]");
		$display("Expect: 115, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 37;
		pixel_array_in[0][2] = 17;
		pixel_array_in[0][3] = 43;
		pixel_array_in[1][0] = 42;
		pixel_array_in[1][1] = 14;
		pixel_array_in[1][2] = 19;
		pixel_array_in[1][3] = 26;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 11;
		pixel_array_in[3][1] = 4;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 38;
		#10;
		
		$display("Input: \n[[17, 16, 23, 57],\n[14, 6, 27, 25],\n[22, 14, 3, 26],\n[40, 55, 29, 32]]");
		$display("Expect: 29, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 3;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 38;
		pixel_array_in[0][3] = 50;
		pixel_array_in[1][0] = 50;
		pixel_array_in[1][1] = 29;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 61;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 33;
		pixel_array_in[3][2] = 5;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[9, 10, 45, 4],\n[42, 4, 35, 30],\n[23, 57, 24, 51],\n[7, 34, 48, 5]]");
		$display("Expect: 120, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 49;
		pixel_array_in[0][1] = 30;
		pixel_array_in[0][2] = 26;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 18;
		pixel_array_in[1][1] = 18;
		pixel_array_in[1][2] = 4;
		pixel_array_in[1][3] = 7;
		pixel_array_in[2][0] = 29;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 29;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 19;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 53;
		#10;
		
		$display("Input: \n[[11, 13, 47, 41],\n[35, 15, 57, 8],\n[60, 27, 54, 40],\n[58, 43, 26, 43]]");
		$display("Expect: 106, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 7;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 10;
		pixel_array_in[0][3] = 21;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 22;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 8;
		#10;
		
		$display("Input: \n[[25, 37, 17, 43],\n[42, 14, 19, 26],\n[30, 23, 17, 30],\n[11, 4, 0, 38]]");
		$display("Expect: 67, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 52;
		pixel_array_in[0][1] = 36;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 24;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 54;
		pixel_array_in[2][2] = 55;
		pixel_array_in[2][3] = 4;
		pixel_array_in[3][0] = 50;
		pixel_array_in[3][1] = 21;
		pixel_array_in[3][2] = 9;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[3, 7, 38, 50],\n[50, 29, 56, 61],\n[1, 45, 7, 9],\n[31, 33, 5, 52]]");
		$display("Expect: 154, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 50;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 18;
		pixel_array_in[0][3] = 27;
		pixel_array_in[1][0] = 52;
		pixel_array_in[1][1] = 43;
		pixel_array_in[1][2] = 34;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 55;
		pixel_array_in[2][1] = 52;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 6;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 8;
		#10;
		
		$display("Input: \n[[49, 30, 26, 15],\n[18, 18, 4, 7],\n[29, 55, 29, 42],\n[38, 19, 56, 53]]");
		$display("Expect: 136, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 6;
		pixel_array_in[0][1] = 9;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 51;
		pixel_array_in[1][2] = 12;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 28;
		pixel_array_in[2][1] = 26;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 55;
		pixel_array_in[3][1] = 51;
		pixel_array_in[3][2] = 43;
		pixel_array_in[3][3] = 28;
		#10;
		
		$display("Input: \n[[7, 0, 10, 21],\n[13, 37, 25, 6],\n[43, 22, 49, 62],\n[38, 48, 59, 8]]");
		$display("Expect: 127, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 24;
		pixel_array_in[0][2] = 54;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 14;
		pixel_array_in[1][1] = 17;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 16;
		pixel_array_in[2][0] = 54;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 46;
		pixel_array_in[2][3] = 13;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 2;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 28;
		#10;
		
		$display("Input: \n[[52, 36, 55, 42],\n[38, 1, 24, 46],\n[50, 54, 55, 4],\n[50, 21, 9, 44]]");
		$display("Expect: 117, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 6;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 31;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 23;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 53;
		pixel_array_in[1][3] = 10;
		pixel_array_in[2][0] = 4;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 4;
		pixel_array_in[3][1] = 33;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 59;
		#10;
		
		$display("Input: \n[[50, 10, 18, 27],\n[52, 43, 34, 6],\n[55, 52, 62, 6],\n[41, 26, 42, 8]]");
		$display("Expect: 207, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 30;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 60;
		pixel_array_in[0][3] = 46;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 19;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 25;
		pixel_array_in[2][1] = 27;
		pixel_array_in[2][2] = 1;
		pixel_array_in[2][3] = 40;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 20;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[6, 9, 13, 57],\n[38, 51, 12, 15],\n[28, 26, 52, 42],\n[55, 51, 43, 28]]");
		$display("Expect: 154, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 60;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 28;
		pixel_array_in[1][0] = 62;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 7;
		pixel_array_in[2][1] = 4;
		pixel_array_in[2][2] = 13;
		pixel_array_in[2][3] = 11;
		pixel_array_in[3][0] = 55;
		pixel_array_in[3][1] = 39;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[22, 24, 54, 8],\n[14, 17, 0, 16],\n[54, 45, 46, 13],\n[46, 2, 27, 28]]");
		$display("Expect: 123, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 4;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 46;
		pixel_array_in[0][3] = 35;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 7;
		pixel_array_in[1][3] = 61;
		pixel_array_in[2][0] = 17;
		pixel_array_in[2][1] = 14;
		pixel_array_in[2][2] = 29;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 18;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 57;
		pixel_array_in[3][3] = 11;
		#10;
		
		$display("Input: \n[[6, 32, 31, 12],\n[23, 1, 53, 10],\n[4, 40, 19, 44],\n[4, 33, 2, 59]]");
		$display("Expect: 94, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 3;
		pixel_array_in[0][1] = 1;
		pixel_array_in[0][2] = 49;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 43;
		pixel_array_in[1][3] = 53;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 5;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 4;
		pixel_array_in[3][3] = 3;
		#10;
		
		$display("Input: \n[[30, 19, 60, 46],\n[31, 27, 19, 4],\n[25, 27, 1, 40],\n[40, 38, 20, 33]]");
		$display("Expect: 89, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 59;
		pixel_array_in[0][2] = 42;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 15;
		pixel_array_in[1][1] = 56;
		pixel_array_in[1][2] = 38;
		pixel_array_in[1][3] = 5;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 18;
		pixel_array_in[3][3] = 14;
		#10;
		
		$display("Input: \n[[15, 60, 23, 28],\n[62, 50, 30, 4],\n[7, 4, 13, 11],\n[55, 39, 0, 60]]");
		$display("Expect: 94, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 47;
		pixel_array_in[0][2] = 49;
		pixel_array_in[0][3] = 14;
		pixel_array_in[1][0] = 6;
		pixel_array_in[1][1] = 20;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 20;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 33;
		pixel_array_in[2][2] = 56;
		pixel_array_in[2][3] = 7;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 61;
		#10;
		
		$display("Input: \n[[4, 19, 46, 35],\n[9, 54, 7, 61],\n[17, 14, 29, 9],\n[18, 14, 57, 11]]");
		$display("Expect: 131, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 36;
		pixel_array_in[0][1] = 22;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 43;
		pixel_array_in[1][0] = 60;
		pixel_array_in[1][1] = 15;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 50;
		pixel_array_in[2][0] = 62;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 12;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 32;
		#10;
		
		$display("Input: \n[[3, 1, 49, 59],\n[38, 35, 43, 53],\n[24, 57, 23, 5],\n[38, 42, 4, 3]]");
		$display("Expect: 189, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 4;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 3;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 51;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 56;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 62;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[32, 59, 42, 10],\n[15, 56, 38, 5],\n[5, 38, 30, 42],\n[40, 0, 18, 14]]");
		$display("Expect: 197, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 57;
		pixel_array_in[0][3] = 28;
		pixel_array_in[1][0] = 15;
		pixel_array_in[1][1] = 47;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 50;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 19;
		pixel_array_in[2][2] = 29;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 62;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 14;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[9, 47, 49, 14],\n[6, 20, 39, 20],\n[10, 33, 56, 7],\n[38, 34, 55, 61]]");
		$display("Expect: 125, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 47;
		pixel_array_in[0][3] = 56;
		pixel_array_in[1][0] = 56;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 54;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 47;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 14;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[36, 22, 7, 43],\n[60, 15, 0, 50],\n[62, 12, 30, 18],\n[10, 12, 17, 32]]");
		$display("Expect: 37, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 13;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 33;
		pixel_array_in[0][3] = 52;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 3;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 6;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 36;
		pixel_array_in[2][3] = 60;
		pixel_array_in[3][0] = 62;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 5;
		#10;
		
		$display("Input: \n[[4, 56, 34, 8],\n[46, 3, 5, 51],\n[5, 56, 30, 62],\n[61, 62, 32, 2]]");
		$display("Expect: 90, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 48;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 42;
		pixel_array_in[0][3] = 13;
		pixel_array_in[1][0] = 33;
		pixel_array_in[1][1] = 38;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 37;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 54;
		#10;
		
		$display("Input: \n[[8, 17, 57, 28],\n[15, 47, 39, 50],\n[14, 19, 29, 9],\n[62, 50, 14, 39]]");
		$display("Expect: 138, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 17;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 60;
		pixel_array_in[1][0] = 7;
		pixel_array_in[1][1] = 18;
		pixel_array_in[1][2] = 7;
		pixel_array_in[1][3] = 24;
		pixel_array_in[2][0] = 16;
		pixel_array_in[2][1] = 16;
		pixel_array_in[2][2] = 12;
		pixel_array_in[2][3] = 7;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 59;
		#10;
		
		$display("Input: \n[[19, 52, 47, 56],\n[56, 32, 32, 54],\n[50, 47, 17, 14],\n[32, 25, 7, 60]]");
		$display("Expect: 140, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 3;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 13;
		pixel_array_in[1][0] = 59;
		pixel_array_in[1][1] = 22;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 55;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 27;
		pixel_array_in[3][0] = 22;
		pixel_array_in[3][1] = 31;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[13, 17, 33, 52],\n[22, 3, 32, 39],\n[6, 36, 36, 60],\n[62, 45, 61, 5]]");
		$display("Expect: 83, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 9;
		pixel_array_in[0][2] = 26;
		pixel_array_in[0][3] = 13;
		pixel_array_in[1][0] = 19;
		pixel_array_in[1][1] = 58;
		pixel_array_in[1][2] = 58;
		pixel_array_in[1][3] = 7;
		pixel_array_in[2][0] = 55;
		pixel_array_in[2][1] = 50;
		pixel_array_in[2][2] = 55;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 21;
		pixel_array_in[3][3] = 24;
		#10;
		
		$display("Input: \n[[48, 0, 42, 13],\n[33, 38, 36, 29],\n[39, 37, 43, 39],\n[29, 57, 17, 54]]");
		$display("Expect: 157, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 26;
		pixel_array_in[0][1] = 6;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 20;
		pixel_array_in[1][0] = 24;
		pixel_array_in[1][1] = 44;
		pixel_array_in[1][2] = 17;
		pixel_array_in[1][3] = 43;
		pixel_array_in[2][0] = 21;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 2;
		pixel_array_in[3][1] = 8;
		pixel_array_in[3][2] = 62;
		pixel_array_in[3][3] = 48;
		#10;
		
		$display("Input: \n[[17, 10, 55, 60],\n[7, 18, 7, 24],\n[16, 16, 12, 7],\n[23, 14, 51, 59]]");
		$display("Expect: 61, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 43;
		pixel_array_in[0][1] = 24;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 5;
		pixel_array_in[1][0] = 53;
		pixel_array_in[1][1] = 62;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 8;
		pixel_array_in[2][0] = 16;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 14;
		pixel_array_in[2][3] = 22;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 52;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 59;
		#10;
		
		$display("Input: \n[[22, 3, 12, 13],\n[59, 22, 0, 46],\n[55, 23, 61, 27],\n[22, 31, 15, 56]]");
		$display("Expect: 89, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 22;
		pixel_array_in[0][3] = 37;
		pixel_array_in[1][0] = 2;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 31;
		pixel_array_in[2][2] = 31;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 61;
		pixel_array_in[3][2] = 10;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[9, 9, 26, 13],\n[19, 58, 58, 7],\n[55, 50, 55, 18],\n[52, 18, 21, 24]]");
		$display("Expect: 248, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 56;
		pixel_array_in[0][1] = 46;
		pixel_array_in[0][2] = 20;
		pixel_array_in[0][3] = 26;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 26;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 23;
		pixel_array_in[2][0] = 28;
		pixel_array_in[2][1] = 21;
		pixel_array_in[2][2] = 45;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 60;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 37;
		#10;
		
		$display("Input: \n[[26, 6, 51, 20],\n[24, 44, 17, 43],\n[21, 17, 57, 24],\n[2, 8, 62, 48]]");
		$display("Expect: 137, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 20;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 47;
		pixel_array_in[1][2] = 1;
		pixel_array_in[1][3] = 55;
		pixel_array_in[2][0] = 59;
		pixel_array_in[2][1] = 49;
		pixel_array_in[2][2] = 35;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 44;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[43, 24, 21, 5],\n[53, 62, 56, 8],\n[16, 55, 14, 22],\n[29, 52, 6, 59]]");
		$display("Expect: 235, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 5;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 21;
		pixel_array_in[2][0] = 46;
		pixel_array_in[2][1] = 47;
		pixel_array_in[2][2] = 46;
		pixel_array_in[2][3] = 45;
		pixel_array_in[3][0] = 6;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 31;
		pixel_array_in[3][3] = 40;
		#10;
		
		$display("Input: \n[[22, 56, 22, 37],\n[2, 23, 56, 12],\n[30, 31, 31, 49],\n[36, 61, 10, 27]]");
		$display("Expect: 115, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 5;
		pixel_array_in[0][1] = 27;
		pixel_array_in[0][2] = 44;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 40;
		pixel_array_in[1][1] = 5;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 5;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 19;
		pixel_array_in[3][0] = 1;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[56, 46, 20, 26],\n[11, 26, 10, 23],\n[28, 21, 45, 53],\n[60, 37, 7, 37]]");
		$display("Expect: 92, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 42;
		pixel_array_in[0][1] = 3;
		pixel_array_in[0][2] = 11;
		pixel_array_in[0][3] = 26;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 51;
		pixel_array_in[2][1] = 4;
		pixel_array_in[2][2] = 10;
		pixel_array_in[2][3] = 29;
		pixel_array_in[3][0] = 34;
		pixel_array_in[3][1] = 4;
		pixel_array_in[3][2] = 54;
		pixel_array_in[3][3] = 49;
		#10;
		
		$display("Input: \n[[20, 18, 12, 10],\n[11, 47, 1, 55],\n[59, 49, 35, 30],\n[5, 48, 44, 20]]");
		$display("Expect: 173, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 26;
		pixel_array_in[0][1] = 47;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 37;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 24;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 25;
		pixel_array_in[3][3] = 37;
		#10;
		
		$display("Input: \n[[53, 32, 52, 39],\n[5, 7, 32, 21],\n[46, 47, 46, 45],\n[6, 59, 31, 40]]");
		$display("Expect: 110, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 2;
		pixel_array_in[0][2] = 36;
		pixel_array_in[0][3] = 11;
		pixel_array_in[1][0] = 62;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 40;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 34;
		#10;
		
		$display("Input: \n[[5, 27, 44, 12],\n[40, 5, 5, 32],\n[40, 5, 57, 19],\n[1, 18, 60, 39]]");
		$display("Expect: 20, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 20;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 9;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 54;
		pixel_array_in[1][1] = 58;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 29;
		pixel_array_in[2][1] = 20;
		pixel_array_in[2][2] = 20;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 9;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 22;
		#10;
		
		$display("Input: \n[[42, 3, 11, 26],\n[46, 12, 30, 38],\n[51, 4, 10, 29],\n[34, 4, 54, 49]]");
		$display("Expect: 29, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 29;
		pixel_array_in[0][2] = 61;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 62;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 7;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 61;
		pixel_array_in[2][2] = 39;
		pixel_array_in[2][3] = 51;
		pixel_array_in[3][0] = 9;
		pixel_array_in[3][1] = 5;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 46;
		#10;
		
		$display("Input: \n[[26, 47, 7, 58],\n[37, 27, 37, 24],\n[42, 35, 49, 43],\n[17, 37, 25, 37]]");
		$display("Expect: 130, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 35;
		pixel_array_in[0][2] = 38;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 35;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 4;
		pixel_array_in[2][1] = 53;
		pixel_array_in[2][2] = 36;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 34;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 14;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[22, 2, 36, 11],\n[62, 25, 15, 6],\n[10, 12, 17, 40],\n[29, 58, 12, 34]]");
		$display("Expect: 60, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 61;
		pixel_array_in[1][3] = 31;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 13;
		pixel_array_in[2][3] = 21;
		pixel_array_in[3][0] = 59;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 8;
		#10;
		
		$display("Input: \n[[20, 25, 9, 1],\n[54, 58, 50, 56],\n[29, 20, 20, 10],\n[9, 28, 59, 22]]");
		$display("Expect: 156, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 7;
		pixel_array_in[0][1] = 39;
		pixel_array_in[0][2] = 20;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 30;
		pixel_array_in[1][1] = 36;
		pixel_array_in[1][2] = 43;
		pixel_array_in[1][3] = 11;
		pixel_array_in[2][0] = 44;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 38;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 41;
		pixel_array_in[3][3] = 62;
		#10;
		
		$display("Input: \n[[61, 29, 61, 15],\n[62, 45, 56, 7],\n[31, 61, 39, 51],\n[9, 5, 12, 46]]");
		$display("Expect: 227, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 51;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 33;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 36;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 13;
		pixel_array_in[3][0] = 58;
		pixel_array_in[3][1] = 36;
		pixel_array_in[3][2] = 46;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[57, 35, 38, 1],\n[11, 60, 35, 25],\n[4, 53, 36, 49],\n[34, 25, 14, 2]]");
		$display("Expect: 235, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 51;
		pixel_array_in[0][2] = 20;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 34;
		pixel_array_in[1][3] = 31;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 29;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 17;
		pixel_array_in[3][0] = 30;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 22;
		#10;
		
		$display("Input: \n[[22, 54, 23, 2],\n[44, 35, 61, 31],\n[22, 10, 13, 21],\n[59, 14, 3, 8]]");
		$display("Expect: 97, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 56;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 43;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 42;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 1;
		pixel_array_in[2][0] = 41;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 56;
		pixel_array_in[3][0] = 60;
		pixel_array_in[3][1] = 35;
		pixel_array_in[3][2] = 34;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[7, 39, 20, 33],\n[30, 36, 43, 11],\n[44, 44, 0, 38],\n[23, 6, 41, 62]]");
		$display("Expect: 151, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 22;
		pixel_array_in[0][2] = 8;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 22;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 28;
		pixel_array_in[2][2] = 18;
		pixel_array_in[2][3] = 58;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 27;
		pixel_array_in[3][2] = 30;
		pixel_array_in[3][3] = 24;
		#10;
		
		$display("Input: \n[[51, 19, 4, 44],\n[33, 45, 5, 36],\n[12, 17, 47, 13],\n[58, 36, 46, 27]]");
		$display("Expect: 125, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 7;
		pixel_array_in[0][1] = 49;
		pixel_array_in[0][2] = 6;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 53;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 20;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 28;
		pixel_array_in[2][2] = 45;
		pixel_array_in[2][3] = 28;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 1;
		pixel_array_in[3][2] = 38;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[8, 51, 20, 33],\n[38, 54, 34, 31],\n[0, 29, 43, 17],\n[30, 37, 7, 22]]");
		$display("Expect: 172, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 23;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 60;
		pixel_array_in[0][3] = 47;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 18;
		pixel_array_in[1][2] = 9;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 46;
		pixel_array_in[2][1] = 34;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 50;
		pixel_array_in[3][0] = 43;
		pixel_array_in[3][1] = 12;
		pixel_array_in[3][2] = 4;
		pixel_array_in[3][3] = 4;
		#10;
		
		$display("Input: \n[[56, 7, 43, 15],\n[42, 45, 36, 1],\n[41, 45, 0, 56],\n[60, 35, 34, 42]]");
		$display("Expect: 166, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 39;
		pixel_array_in[0][1] = 5;
		pixel_array_in[0][2] = 20;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 15;
		pixel_array_in[1][1] = 57;
		pixel_array_in[1][2] = 52;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 36;
		pixel_array_in[2][1] = 46;
		pixel_array_in[2][2] = 4;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 45;
		pixel_array_in[3][1] = 41;
		pixel_array_in[3][2] = 1;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[22, 22, 8, 2],\n[22, 1, 11, 22],\n[24, 28, 18, 58],\n[10, 27, 30, 24]]");
		$display("Expect: 47, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 49;
		pixel_array_in[0][1] = 8;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 30;
		pixel_array_in[1][0] = 19;
		pixel_array_in[1][1] = 13;
		pixel_array_in[1][2] = 43;
		pixel_array_in[1][3] = 60;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 39;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 10;
		pixel_array_in[3][2] = 1;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[7, 49, 6, 45],\n[53, 23, 15, 20],\n[15, 28, 45, 28],\n[42, 1, 38, 1]]");
		$display("Expect: 104, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 44;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 40;
		pixel_array_in[0][3] = 34;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 23;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 54;
		pixel_array_in[2][1] = 22;
		pixel_array_in[2][2] = 59;
		pixel_array_in[2][3] = 60;
		pixel_array_in[3][0] = 50;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[23, 45, 60, 47],\n[31, 18, 9, 18],\n[46, 34, 57, 50],\n[43, 12, 4, 4]]");
		$display("Expect: 104, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 27;
		pixel_array_in[0][1] = 13;
		pixel_array_in[0][2] = 54;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 41;
		pixel_array_in[1][1] = 10;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 57;
		pixel_array_in[2][0] = 7;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 2;
		pixel_array_in[2][3] = 35;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 22;
		#10;
		
		$display("Input: \n[[39, 5, 20, 44],\n[15, 57, 52, 6],\n[36, 46, 4, 43],\n[45, 41, 1, 58]]");
		$display("Expect: 209, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 54;
		pixel_array_in[0][1] = 11;
		pixel_array_in[0][2] = 9;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 24;
		pixel_array_in[1][1] = 62;
		pixel_array_in[1][2] = 51;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 13;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 34;
		pixel_array_in[2][3] = 5;
		pixel_array_in[3][0] = 47;
		pixel_array_in[3][1] = 4;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 19;
		#10;
		
		$display("Input: \n[[49, 8, 51, 30],\n[19, 13, 43, 60],\n[42, 12, 39, 25],\n[42, 10, 1, 7]]");
		$display("Expect: 71, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 12;
		pixel_array_in[0][1] = 39;
		pixel_array_in[0][2] = 37;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 17;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 60;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 62;
		pixel_array_in[2][2] = 10;
		pixel_array_in[2][3] = 21;
		pixel_array_in[3][0] = 47;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 37;
		pixel_array_in[3][3] = 50;
		#10;
		
		$display("Input: \n[[44, 28, 40, 34],\n[31, 33, 23, 62],\n[54, 22, 59, 60],\n[50, 26, 42, 1]]");
		$display("Expect: 114, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 58;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 37;
		pixel_array_in[0][3] = 47;
		pixel_array_in[1][0] = 51;
		pixel_array_in[1][1] = 17;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 56;
		pixel_array_in[2][1] = 6;
		pixel_array_in[2][2] = 60;
		pixel_array_in[2][3] = 47;
		pixel_array_in[3][0] = 8;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 49;
		#10;
		
		$display("Input: \n[[27, 13, 54, 25],\n[41, 10, 30, 57],\n[7, 12, 2, 35],\n[61, 26, 55, 22]]");
		$display("Expect: 33, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 4;
		pixel_array_in[0][1] = 4;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 41;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 48;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 28;
		pixel_array_in[2][1] = 27;
		pixel_array_in[2][2] = 10;
		pixel_array_in[2][3] = 15;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 11;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 59;
		#10;
		
		$display("Input: \n[[54, 11, 9, 45],\n[24, 62, 51, 56],\n[13, 32, 34, 5],\n[47, 4, 42, 19]]");
		$display("Expect: 213, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 31;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 14;
		pixel_array_in[1][2] = 58;
		pixel_array_in[1][3] = 59;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 26;
		pixel_array_in[2][2] = 37;
		pixel_array_in[2][3] = 2;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 32;
		#10;
		
		$display("Input: \n[[12, 39, 37, 33],\n[17, 7, 30, 60],\n[22, 62, 10, 21],\n[47, 32, 37, 50]]");
		$display("Expect: 126, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 48;
		pixel_array_in[0][1] = 13;
		pixel_array_in[0][2] = 53;
		pixel_array_in[0][3] = 3;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 60;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 61;
		pixel_array_in[2][1] = 27;
		pixel_array_in[2][2] = 2;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 41;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[58, 7, 37, 47],\n[51, 17, 11, 62],\n[56, 6, 60, 47],\n[8, 26, 27, 49]]");
		$display("Expect: 49, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 52;
		pixel_array_in[0][1] = 34;
		pixel_array_in[0][2] = 11;
		pixel_array_in[0][3] = 29;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 3;
		pixel_array_in[2][0] = 9;
		pixel_array_in[2][1] = 60;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 45;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 62;
		pixel_array_in[3][3] = 30;
		#10;
		
		$display("Input: \n[[4, 4, 51, 41],\n[41, 0, 48, 46],\n[28, 27, 10, 15],\n[19, 11, 36, 59]]");
		$display("Expect: 61, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 34;
		pixel_array_in[0][1] = 62;
		pixel_array_in[0][2] = 25;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 55;
		pixel_array_in[1][2] = 61;
		pixel_array_in[1][3] = 20;
		pixel_array_in[2][0] = 52;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 12;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 61;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[29, 10, 4, 31],\n[38, 14, 58, 59],\n[60, 26, 37, 2],\n[29, 0, 36, 32]]");
		$display("Expect: 104, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 40;
		pixel_array_in[0][1] = 12;
		pixel_array_in[0][2] = 3;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 60;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 33;
		pixel_array_in[2][0] = 61;
		pixel_array_in[2][1] = 5;
		pixel_array_in[2][2] = 16;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 21;
		pixel_array_in[3][1] = 51;
		pixel_array_in[3][2] = 52;
		pixel_array_in[3][3] = 24;
		#10;
		
		$display("Input: \n[[48, 13, 53, 3],\n[13, 45, 60, 39],\n[61, 27, 2, 41],\n[32, 38, 41, 58]]");
		$display("Expect: 141, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 33;
		pixel_array_in[0][1] = 50;
		pixel_array_in[0][2] = 44;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 48;
		pixel_array_in[1][1] = 42;
		pixel_array_in[1][2] = 49;
		pixel_array_in[1][3] = 28;
		pixel_array_in[2][0] = 46;
		pixel_array_in[2][1] = 14;
		pixel_array_in[2][2] = 38;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[52, 34, 11, 29],\n[61, 25, 37, 3],\n[9, 60, 49, 53],\n[45, 18, 62, 30]]");
		$display("Expect: 182, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 5;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 21;
		pixel_array_in[1][3] = 22;
		pixel_array_in[2][0] = 41;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 58;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 37;
		#10;
		
		$display("Input: \n[[34, 62, 25, 41],\n[28, 55, 61, 20],\n[52, 11, 17, 12],\n[17, 61, 55, 16]]");
		$display("Expect: 124, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 13;
		pixel_array_in[0][1] = 14;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 21;
		pixel_array_in[1][1] = 47;
		pixel_array_in[1][2] = 43;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 44;
		pixel_array_in[2][1] = 51;
		pixel_array_in[2][2] = 21;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 47;
		pixel_array_in[3][3] = 36;
		#10;
		
		$display("Input: \n[[40, 12, 3, 2],\n[60, 54, 13, 33],\n[61, 5, 16, 41],\n[21, 51, 52, 24]]");
		$display("Expect: 91, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 2;
		pixel_array_in[0][1] = 22;
		pixel_array_in[0][2] = 25;
		pixel_array_in[0][3] = 27;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 47;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 53;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 19;
		pixel_array_in[2][2] = 26;
		pixel_array_in[2][3] = 34;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 27;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 22;
		#10;
		
		$display("Input: \n[[33, 50, 44, 55],\n[48, 42, 49, 28],\n[46, 14, 38, 32],\n[13, 50, 55, 27]]");
		$display("Expect: 109, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 31;
		pixel_array_in[0][1] = 30;
		pixel_array_in[0][2] = 61;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 39;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 44;
		pixel_array_in[2][1] = 43;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 54;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[25, 5, 13, 12],\n[32, 7, 21, 22],\n[41, 45, 47, 58],\n[23, 13, 12, 37]]");
		$display("Expect: 116, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 45;
		pixel_array_in[0][1] = 35;
		pixel_array_in[0][2] = 41;
		pixel_array_in[0][3] = 23;
		pixel_array_in[1][0] = 7;
		pixel_array_in[1][1] = 30;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 3;
		pixel_array_in[2][0] = 19;
		pixel_array_in[2][1] = 29;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 57;
		pixel_array_in[3][1] = 49;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 46;
		#10;
		
		$display("Input: \n[[13, 14, 19, 40],\n[21, 47, 43, 25],\n[44, 51, 21, 42],\n[40, 28, 47, 36]]");
		$display("Expect: 198, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 54;
		pixel_array_in[0][1] = 33;
		pixel_array_in[0][2] = 50;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 46;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 6;
		pixel_array_in[2][1] = 47;
		pixel_array_in[2][2] = 53;
		pixel_array_in[2][3] = 23;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 31;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[2, 22, 25, 27],\n[31, 47, 30, 53],\n[24, 19, 26, 34],\n[46, 27, 32, 22]]");
		$display("Expect: 131, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 36;
		pixel_array_in[0][1] = 62;
		pixel_array_in[0][2] = 40;
		pixel_array_in[0][3] = 24;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 31;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 33;
		pixel_array_in[2][0] = 2;
		pixel_array_in[2][1] = 31;
		pixel_array_in[2][2] = 45;
		pixel_array_in[2][3] = 29;
		pixel_array_in[3][0] = 24;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 15;
		#10;
		
		$display("Input: \n[[31, 30, 61, 53],\n[39, 12, 50, 44],\n[44, 43, 43, 43],\n[54, 14, 2, 44]]");
		$display("Expect: 125, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 17;
		pixel_array_in[0][1] = 44;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 4;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 1;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 23;
		pixel_array_in[2][1] = 48;
		pixel_array_in[2][2] = 3;
		pixel_array_in[2][3] = 61;
		pixel_array_in[3][0] = 33;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 43;
		#10;
		
		$display("Input: \n[[45, 35, 41, 23],\n[7, 30, 39, 3],\n[19, 29, 57, 49],\n[57, 49, 48, 46]]");
		$display("Expect: 135, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 45;
		pixel_array_in[1][1] = 34;
		pixel_array_in[1][2] = 49;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 52;
		pixel_array_in[2][1] = 39;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 22;
		pixel_array_in[3][0] = 22;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[54, 33, 50, 18],\n[11, 46, 3, 18],\n[6, 47, 53, 23],\n[10, 57, 31, 7]]");
		$display("Expect: 182, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 1;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 36;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 17;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 18;
		#10;
		
		$display("Input: \n[[36, 62, 40, 24],\n[61, 31, 10, 33],\n[2, 31, 45, 29],\n[24, 28, 36, 15]]");
		$display("Expect: 113, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 45;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 28;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 30;
		pixel_array_in[1][1] = 34;
		pixel_array_in[1][2] = 57;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[17, 44, 52, 2],\n[4, 54, 1, 18],\n[23, 48, 3, 61],\n[33, 26, 0, 43]]");
		$display("Expect: 175, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 38;
		pixel_array_in[0][1] = 9;
		pixel_array_in[0][2] = 37;
		pixel_array_in[0][3] = 49;
		pixel_array_in[1][0] = 55;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 45;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 18;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 10;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[53, 7, 13, 40],\n[45, 34, 49, 48],\n[52, 39, 43, 22],\n[22, 58, 60, 42]]");
		$display("Expect: 153, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 2;
		pixel_array_in[0][1] = 44;
		pixel_array_in[0][2] = 5;
		pixel_array_in[0][3] = 28;
		pixel_array_in[1][0] = 52;
		pixel_array_in[1][1] = 24;
		pixel_array_in[1][2] = 14;
		pixel_array_in[1][3] = 45;
		pixel_array_in[2][0] = 32;
		pixel_array_in[2][1] = 58;
		pixel_array_in[2][2] = 40;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 17;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[19, 58, 21, 41],\n[47, 33, 1, 12],\n[36, 10, 19, 17],\n[32, 30, 48, 18]]");
		$display("Expect: 57, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 35;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 58;
		pixel_array_in[0][3] = 37;
		pixel_array_in[1][0] = 16;
		pixel_array_in[1][1] = 10;
		pixel_array_in[1][2] = 24;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 55;
		pixel_array_in[2][1] = 21;
		pixel_array_in[2][2] = 45;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 54;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 1;
		pixel_array_in[3][3] = 10;
		#10;
		
		$display("Input: \n[[45, 45, 28, 58],\n[30, 34, 57, 15],\n[0, 40, 30, 10],\n[38, 57, 42, 52]]");
		$display("Expect: 158, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 54;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 60;
		pixel_array_in[1][1] = 47;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 48;
		pixel_array_in[2][1] = 14;
		pixel_array_in[2][2] = 37;
		pixel_array_in[2][3] = 12;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 51;
		#10;
		
		$display("Input: \n[[38, 9, 37, 49],\n[55, 37, 5, 62],\n[45, 13, 18, 9],\n[13, 10, 29, 35]]");
		$display("Expect: 83, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 62;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 61;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 30;
		pixel_array_in[1][1] = 15;
		pixel_array_in[1][2] = 26;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 37;
		pixel_array_in[2][1] = 27;
		pixel_array_in[2][2] = 11;
		pixel_array_in[2][3] = 56;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 43;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 22;
		#10;
		
		$display("Input: \n[[2, 44, 5, 28],\n[52, 24, 14, 45],\n[32, 58, 40, 25],\n[61, 17, 17, 2]]");
		$display("Expect: 157, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 48;
		pixel_array_in[0][1] = 57;
		pixel_array_in[0][2] = 38;
		pixel_array_in[0][3] = 32;
		pixel_array_in[1][0] = 59;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 34;
		pixel_array_in[3][1] = 29;
		pixel_array_in[3][2] = 8;
		pixel_array_in[3][3] = 55;
		#10;
		
		$display("Input: \n[[35, 26, 58, 37],\n[16, 10, 24, 47],\n[55, 21, 45, 39],\n[54, 55, 1, 10]]");
		$display("Expect: 60, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 12;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 53;
		pixel_array_in[1][1] = 5;
		pixel_array_in[1][2] = 24;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 8;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 14;
		pixel_array_in[2][3] = 26;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 54;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 13;
		#10;
		
		$display("Input: \n[[19, 28, 54, 53],\n[60, 47, 3, 17],\n[48, 14, 37, 12],\n[13, 37, 2, 51]]");
		$display("Expect: 105, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 54;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 11;
		pixel_array_in[1][0] = 20;
		pixel_array_in[1][1] = 16;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 28;
		pixel_array_in[2][0] = 35;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 50;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 22;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[62, 10, 61, 8],\n[30, 15, 26, 38],\n[37, 27, 11, 56],\n[29, 43, 12, 22]]");
		$display("Expect: 71, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 47;
		pixel_array_in[0][2] = 10;
		pixel_array_in[0][3] = 50;
		pixel_array_in[1][0] = 36;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 23;
		pixel_array_in[1][3] = 20;
		pixel_array_in[2][0] = 37;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 25;
		pixel_array_in[2][3] = 27;
		pixel_array_in[3][0] = 18;
		pixel_array_in[3][1] = 1;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[48, 57, 38, 32],\n[59, 49, 22, 39],\n[22, 40, 43, 30],\n[34, 29, 8, 55]]");
		$display("Expect: 171, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 42;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 9;
		pixel_array_in[1][2] = 52;
		pixel_array_in[1][3] = 9;
		pixel_array_in[2][0] = 58;
		pixel_array_in[2][1] = 39;
		pixel_array_in[2][2] = 28;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 21;
		pixel_array_in[3][2] = 40;
		pixel_array_in[3][3] = 55;
		#10;
		
		$display("Input: \n[[12, 56, 55, 39],\n[53, 5, 24, 48],\n[8, 57, 14, 26],\n[46, 54, 45, 13]]");
		$display("Expect: 98, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 20;
		pixel_array_in[0][1] = 14;
		pixel_array_in[0][2] = 49;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 53;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 36;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 53;
		pixel_array_in[2][3] = 11;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 47;
		#10;
		
		$display("Input: \n[[54, 48, 48, 11],\n[20, 16, 5, 28],\n[35, 0, 62, 36],\n[50, 42, 22, 7]]");
		$display("Expect: 31, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 35;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 16;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 2;
		pixel_array_in[2][3] = 6;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 17;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[9, 47, 10, 50],\n[36, 37, 23, 20],\n[37, 57, 25, 27],\n[18, 1, 7, 58]]");
		$display("Expect: 183, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 45;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 38;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 58;
		pixel_array_in[1][3] = 23;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 50;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 23;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 22;
		pixel_array_in[3][2] = 31;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[0, 45, 42, 42],\n[10, 9, 52, 9],\n[58, 39, 28, 41],\n[15, 21, 40, 55]]");
		$display("Expect: 103, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 24;
		pixel_array_in[0][1] = 57;
		pixel_array_in[0][2] = 11;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 12;
		pixel_array_in[1][1] = 38;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 43;
		pixel_array_in[2][0] = 55;
		pixel_array_in[2][1] = 62;
		pixel_array_in[2][2] = 8;
		pixel_array_in[2][3] = 52;
		pixel_array_in[3][0] = 24;
		pixel_array_in[3][1] = 36;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 4;
		#10;
		
		$display("Input: \n[[20, 14, 49, 40],\n[53, 45, 11, 36],\n[12, 35, 53, 11],\n[25, 38, 32, 47]]");
		$display("Expect: 161, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 10;
		pixel_array_in[0][1] = 1;
		pixel_array_in[0][2] = 24;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 25;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 35;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 18;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 17;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[25, 45, 35, 12],\n[28, 16, 32, 56],\n[40, 57, 2, 6],\n[19, 17, 6, 2]]");
		$display("Expect: 130, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 51;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 22;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 56;
		pixel_array_in[1][2] = 20;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 23;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 30;
		#10;
		
		$display("Input: \n[[45, 18, 30, 38],\n[22, 52, 58, 23],\n[12, 50, 54, 23],\n[5, 22, 31, 7]]");
		$display("Expect: 237, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[24, 57, 11, 1],\n[12, 38, 33, 43],\n[55, 62, 8, 52],\n[24, 36, 17, 4]]");
		$display("Expect: 179, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[10, 1, 24, 44],\n[25, 7, 35, 4],\n[43, 18, 62, 25],\n[40, 17, 15, 56]]");
		$display("Expect: 81, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[51, 25, 22, 19],\n[58, 56, 20, 18],\n[50, 38, 5, 9],\n[23, 23, 42, 30]]");
		$display("Expect: 165, Result: %d", pixel_out);
		$display("");
		#10;
		
		
		$display("Finishing Sim"); //print nice message
		$finish;
		
    end
endmodule //counter_tb

`default_nettype wire