`timescale 1ns / 1ps
`default_nettype none

module kernel_5_tb;

    //make logics for inputs and outputs!
    logic clk_in;
    logic rst_in;
    logic valid_in;
    logic [5:0] pixel_array_in [3:0][3:0];
    logic [8:0] pixel_out;

    kernel_5 uut (
        .clk_in(clk_in),
        .p(pixel_array_in),
        .pixel_out(pixel_out)
    );
    always begin
        #5;  //every 5 ns switch...so period of clock is 10 ns...100 MHz clock
        clk_in = !clk_in;
    end

    //initial block...this is our test simulation
    initial begin

		$dumpfile("test/kernel_5.vcd"); //file to store value change dump (vcd)
		$dumpvars(0,kernel_5_tb); //store everything at the current level and below
		$display("Starting Sim"); //print nice message
		clk_in = 0; //initialize clk (super important)
		rst_in = 0; //initialize rst (super important)
		
		#10;  //wait a little bit of time at beginning
		rst_in = 1; //reset system
		#10; //hold high for a few clock cycles
		rst_in=0;
		
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 0;
		#10;
		
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 32;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 32;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 32;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 32;
		#10;
		
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 63;
		#10;
		
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 63;
		#10;
		
		$display("Input: \n[[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0]]");
		$display("Expect: 0, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Input: \n[[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32]]");
		$display("Expect: 128, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 23;
		pixel_array_in[0][1] = 36;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 48;
		pixel_array_in[1][1] = 36;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 37;
		pixel_array_in[2][1] = 30;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 22;
		pixel_array_in[3][3] = 51;
		#10;
		
		$display("Input: \n[[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63]]");
		$display("Expect: 252, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 18;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 26;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 59;
		pixel_array_in[2][1] = 54;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 13;
		pixel_array_in[3][0] = 3;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 26;
		pixel_array_in[3][3] = 21;
		#10;
		
		$display("Input: \n[[63, 0, 0, 63],\n[0, 63, 63, 0],\n[0, 63, 63, 0],\n[63, 0, 0, 63]]");
		$display("Expect: 384>val>255, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 42;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 28;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 25;
		pixel_array_in[1][1] = 20;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 23;
		pixel_array_in[2][0] = 23;
		pixel_array_in[2][1] = 50;
		pixel_array_in[2][2] = 6;
		pixel_array_in[2][3] = 6;
		pixel_array_in[3][0] = 39;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 21;
		pixel_array_in[3][3] = 55;
		#10;
		
		$display("Input: \n[[0, 63, 63, 0],\n[63, 0, 0, 63],\n[63, 0, 0, 63],\n[0, 63, 63, 0]]");
		$display("Expect: val>383, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 13;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 62;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 60;
		pixel_array_in[2][3] = 2;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 51;
		pixel_array_in[3][2] = 40;
		pixel_array_in[3][3] = 30;
		#10;
		
		$display("Input: \n[[23, 36, 14, 39],\n[48, 36, 22, 35],\n[37, 30, 30, 1],\n[17, 13, 22, 51]]");
		$display("Expect: 122, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 28;
		pixel_array_in[0][1] = 47;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 16;
		pixel_array_in[1][0] = 4;
		pixel_array_in[1][1] = 43;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 45;
		pixel_array_in[2][1] = 26;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 48;
		pixel_array_in[3][1] = 15;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[18, 54, 12, 26],\n[38, 25, 10, 29],\n[59, 54, 61, 13],\n[3, 30, 26, 21]]");
		$display("Expect: 154, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 48;
		pixel_array_in[0][1] = 51;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 38;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 37;
		pixel_array_in[2][1] = 9;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 25;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[42, 19, 28, 44],\n[25, 20, 11, 23],\n[23, 50, 6, 6],\n[39, 44, 21, 55]]");
		$display("Expect: 86, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 14;
		pixel_array_in[0][1] = 46;
		pixel_array_in[0][2] = 10;
		pixel_array_in[0][3] = 24;
		pixel_array_in[1][0] = 40;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 20;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 9;
		pixel_array_in[2][2] = 59;
		pixel_array_in[2][3] = 2;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 10;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[13, 48, 4, 55],\n[61, 62, 50, 56],\n[39, 7, 60, 2],\n[10, 51, 40, 30]]");
		$display("Expect: 185, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 47;
		pixel_array_in[0][2] = 2;
		pixel_array_in[0][3] = 6;
		pixel_array_in[1][0] = 33;
		pixel_array_in[1][1] = 31;
		pixel_array_in[1][2] = 21;
		pixel_array_in[1][3] = 57;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 21;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 20;
		pixel_array_in[3][0] = 7;
		pixel_array_in[3][1] = 33;
		pixel_array_in[3][2] = 10;
		pixel_array_in[3][3] = 49;
		#10;
		
		$display("Input: \n[[28, 47, 19, 16],\n[4, 43, 50, 35],\n[45, 26, 62, 1],\n[48, 15, 36, 12]]");
		$display("Expect: 202, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 11;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 53;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 19;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 19;
		pixel_array_in[2][0] = 8;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 28;
		pixel_array_in[2][3] = 6;
		pixel_array_in[3][0] = 54;
		pixel_array_in[3][1] = 36;
		pixel_array_in[3][2] = 35;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[48, 51, 7, 38],\n[9, 49, 32, 12],\n[37, 9, 22, 62],\n[42, 0, 25, 56]]");
		$display("Expect: 116, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 25;
		pixel_array_in[0][3] = 46;
		pixel_array_in[1][0] = 55;
		pixel_array_in[1][1] = 29;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 2;
		pixel_array_in[2][0] = 18;
		pixel_array_in[2][1] = 16;
		pixel_array_in[2][2] = 40;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 23;
		pixel_array_in[3][2] = 16;
		pixel_array_in[3][3] = 28;
		#10;
		
		$display("Input: \n[[14, 46, 10, 24],\n[40, 28, 20, 62],\n[39, 9, 59, 2],\n[19, 10, 45, 39]]");
		$display("Expect: 112, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 45;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 28;
		pixel_array_in[1][0] = 42;
		pixel_array_in[1][1] = 21;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 47;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 11;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 52;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 57;
		#10;
		
		$display("Input: \n[[25, 47, 2, 6],\n[33, 31, 21, 57],\n[50, 21, 44, 20],\n[7, 33, 10, 49]]");
		$display("Expect: 114, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 33;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 56;
		pixel_array_in[1][1] = 53;
		pixel_array_in[1][2] = 35;
		pixel_array_in[1][3] = 49;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 56;
		pixel_array_in[2][2] = 59;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 52;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[11, 19, 53, 33],\n[19, 60, 10, 19],\n[8, 32, 28, 6],\n[54, 36, 35, 16]]");
		$display("Expect: 138, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 5;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 24;
		pixel_array_in[1][0] = 62;
		pixel_array_in[1][1] = 58;
		pixel_array_in[1][2] = 35;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 45;
		pixel_array_in[2][1] = 39;
		pixel_array_in[2][2] = 48;
		pixel_array_in[2][3] = 19;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 28;
		pixel_array_in[3][3] = 21;
		#10;
		
		$display("Input: \n[[29, 19, 25, 46],\n[55, 29, 30, 2],\n[18, 16, 40, 0],\n[31, 23, 16, 28]]");
		$display("Expect: 125, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 4;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 30;
		pixel_array_in[1][0] = 37;
		pixel_array_in[1][1] = 59;
		pixel_array_in[1][2] = 43;
		pixel_array_in[1][3] = 51;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 49;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 48;
		pixel_array_in[3][0] = 28;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 25;
		#10;
		
		$display("Input: \n[[45, 26, 34, 28],\n[42, 21, 33, 48],\n[5, 47, 22, 11],\n[31, 52, 42, 57]]");
		$display("Expect: 121, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 8;
		pixel_array_in[0][3] = 3;
		pixel_array_in[1][0] = 26;
		pixel_array_in[1][1] = 62;
		pixel_array_in[1][2] = 46;
		pixel_array_in[1][3] = 2;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 24;
		pixel_array_in[2][2] = 20;
		pixel_array_in[2][3] = 50;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 4;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 36;
		#10;
		
		$display("Input: \n[[1, 33, 30, 55],\n[56, 53, 35, 49],\n[12, 56, 59, 53],\n[13, 6, 52, 33]]");
		$display("Expect: 217, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 50;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 31;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 5;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 4;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 49;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 28;
		pixel_array_in[2][3] = 27;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 3;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[5, 56, 0, 24],\n[62, 58, 35, 46],\n[45, 39, 48, 19],\n[17, 42, 28, 21]]");
		$display("Expect: 186, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 5;
		pixel_array_in[0][1] = 42;
		pixel_array_in[0][2] = 20;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 9;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 37;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 1;
		pixel_array_in[3][1] = 24;
		pixel_array_in[3][2] = 62;
		pixel_array_in[3][3] = 10;
		#10;
		
		$display("Input: \n[[8, 4, 34, 30],\n[37, 59, 43, 51],\n[57, 49, 42, 48],\n[28, 38, 48, 25]]");
		$display("Expect: 201, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 4;
		pixel_array_in[0][2] = 44;
		pixel_array_in[0][3] = 5;
		pixel_array_in[1][0] = 15;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 46;
		pixel_array_in[1][3] = 10;
		pixel_array_in[2][0] = 25;
		pixel_array_in[2][1] = 49;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 14;
		pixel_array_in[3][0] = 2;
		pixel_array_in[3][1] = 56;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 3;
		#10;
		
		$display("Input: \n[[29, 10, 8, 3],\n[26, 62, 46, 2],\n[60, 24, 20, 50],\n[31, 4, 56, 36]]");
		$display("Expect: 163, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 24;
		pixel_array_in[0][1] = 46;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 36;
		pixel_array_in[1][2] = 23;
		pixel_array_in[1][3] = 10;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 41;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 20;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 49;
		pixel_array_in[3][3] = 50;
		#10;
		
		$display("Input: \n[[50, 18, 31, 40],\n[5, 54, 4, 62],\n[49, 17, 28, 27],\n[10, 3, 59, 42]]");
		$display("Expect: 96, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 11;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 29;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 53;
		pixel_array_in[1][2] = 38;
		pixel_array_in[1][3] = 51;
		pixel_array_in[2][0] = 35;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 40;
		pixel_array_in[2][3] = 46;
		pixel_array_in[3][0] = 18;
		pixel_array_in[3][1] = 43;
		pixel_array_in[3][2] = 13;
		pixel_array_in[3][3] = 18;
		#10;
		
		$display("Input: \n[[5, 42, 20, 44],\n[57, 45, 9, 18],\n[40, 37, 17, 36],\n[1, 24, 62, 10]]");
		$display("Expect: 95, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 33;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 11;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 17;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 40;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 20;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 21;
		pixel_array_in[3][3] = 21;
		#10;
		
		$display("Input: \n[[19, 4, 44, 5],\n[15, 60, 46, 10],\n[25, 49, 62, 14],\n[2, 56, 12, 3]]");
		$display("Expect: 249, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 27;
		pixel_array_in[0][1] = 44;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 35;
		pixel_array_in[1][1] = 39;
		pixel_array_in[1][2] = 16;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 24;
		pixel_array_in[2][3] = 7;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[24, 46, 21, 8],\n[0, 36, 23, 10],\n[14, 41, 49, 9],\n[20, 30, 49, 50]]");
		$display("Expect: 165, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 31;
		pixel_array_in[0][1] = 50;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 58;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 1;
		pixel_array_in[2][0] = 2;
		pixel_array_in[2][1] = 5;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 45;
		pixel_array_in[3][1] = 4;
		pixel_array_in[3][2] = 41;
		pixel_array_in[3][3] = 34;
		#10;
		
		$display("Input: \n[[8, 11, 45, 29],\n[9, 53, 38, 51],\n[35, 17, 40, 46],\n[18, 43, 13, 18]]");
		$display("Expect: 152, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 47;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 15;
		pixel_array_in[1][1] = 10;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 2;
		pixel_array_in[2][0] = 7;
		pixel_array_in[2][1] = 61;
		pixel_array_in[2][2] = 41;
		pixel_array_in[2][3] = 15;
		pixel_array_in[3][0] = 47;
		pixel_array_in[3][1] = 4;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 32;
		#10;
		
		$display("Input: \n[[33, 17, 52, 36],\n[28, 11, 15, 12],\n[17, 55, 40, 49],\n[20, 55, 21, 21]]");
		$display("Expect: 119, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 62;
		pixel_array_in[0][1] = 6;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 17;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 61;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 8;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 6;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 22;
		pixel_array_in[3][2] = 43;
		pixel_array_in[3][3] = 49;
		#10;
		
		$display("Input: \n[[27, 44, 19, 25],\n[35, 39, 16, 17],\n[5, 13, 24, 7],\n[38, 32, 11, 2]]");
		$display("Expect: 93, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 17;
		pixel_array_in[0][1] = 41;
		pixel_array_in[0][2] = 59;
		pixel_array_in[0][3] = 16;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 40;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 56;
		pixel_array_in[3][0] = 51;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 19;
		pixel_array_in[3][3] = 32;
		#10;
		
		$display("Input: \n[[31, 50, 30, 57],\n[61, 58, 22, 1],\n[2, 5, 42, 44],\n[45, 4, 41, 34]]");
		$display("Expect: 130, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 3;
		pixel_array_in[0][1] = 8;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 20;
		pixel_array_in[1][0] = 39;
		pixel_array_in[1][1] = 4;
		pixel_array_in[1][2] = 42;
		pixel_array_in[1][3] = 30;
		pixel_array_in[2][0] = 18;
		pixel_array_in[2][1] = 43;
		pixel_array_in[2][2] = 21;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 53;
		pixel_array_in[3][1] = 39;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[8, 47, 12, 36],\n[15, 10, 15, 2],\n[7, 61, 41, 15],\n[47, 4, 60, 32]]");
		$display("Expect: 139, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 36;
		pixel_array_in[1][2] = 38;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 53;
		pixel_array_in[2][1] = 22;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 8;
		#10;
		
		$display("Input: \n[[62, 6, 48, 17],\n[10, 61, 15, 8],\n[5, 36, 6, 3],\n[52, 22, 43, 49]]");
		$display("Expect: 131, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 59;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 25;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 37;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 47;
		pixel_array_in[1][3] = 20;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 20;
		pixel_array_in[2][2] = 45;
		pixel_array_in[2][3] = 28;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 50;
		pixel_array_in[3][3] = 36;
		#10;
		
		$display("Input: \n[[17, 41, 59, 16],\n[11, 40, 32, 62],\n[39, 0, 61, 56],\n[51, 25, 19, 32]]");
		$display("Expect: 126, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 49;
		pixel_array_in[0][1] = 3;
		pixel_array_in[0][2] = 39;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 5;
		pixel_array_in[1][1] = 18;
		pixel_array_in[1][2] = 29;
		pixel_array_in[1][3] = 10;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 22;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 62;
		pixel_array_in[3][2] = 16;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[3, 8, 23, 20],\n[39, 4, 42, 30],\n[18, 43, 21, 3],\n[53, 39, 59, 20]]");
		$display("Expect: 109, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 38;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 8;
		pixel_array_in[1][2] = 12;
		pixel_array_in[1][3] = 13;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 34;
		pixel_array_in[3][0] = 7;
		pixel_array_in[3][1] = 20;
		pixel_array_in[3][2] = 53;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[9, 45, 30, 44],\n[10, 36, 38, 0],\n[53, 22, 61, 24],\n[23, 0, 12, 8]]");
		$display("Expect: 175, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 12;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 34;
		pixel_array_in[1][2] = 48;
		pixel_array_in[1][3] = 42;
		pixel_array_in[2][0] = 25;
		pixel_array_in[2][1] = 56;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 48;
		pixel_array_in[3][0] = 6;
		pixel_array_in[3][1] = 49;
		pixel_array_in[3][2] = 1;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[59, 17, 25, 33],\n[37, 54, 47, 20],\n[30, 20, 45, 28],\n[15, 13, 50, 36]]");
		$display("Expect: 181, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 3;
		pixel_array_in[0][1] = 59;
		pixel_array_in[0][2] = 36;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 36;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 30;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 56;
		pixel_array_in[2][2] = 55;
		pixel_array_in[2][3] = 34;
		pixel_array_in[3][0] = 37;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 43;
		#10;
		
		$display("Input: \n[[49, 3, 39, 19],\n[5, 18, 29, 10],\n[50, 22, 49, 43],\n[17, 62, 16, 44]]");
		$display("Expect: 119, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 56;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 42;
		pixel_array_in[1][3] = 58;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 4;
		pixel_array_in[2][2] = 20;
		pixel_array_in[2][3] = 38;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 27;
		pixel_array_in[3][2] = 1;
		pixel_array_in[3][3] = 23;
		#10;
		
		$display("Input: \n[[53, 52, 52, 38],\n[44, 8, 12, 13],\n[57, 57, 22, 34],\n[7, 20, 53, 27]]");
		$display("Expect: 81, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 12;
		pixel_array_in[0][1] = 20;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 18;
		pixel_array_in[1][1] = 58;
		pixel_array_in[1][2] = 41;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 49;
		pixel_array_in[2][1] = 42;
		pixel_array_in[2][2] = 15;
		pixel_array_in[2][3] = 2;
		pixel_array_in[3][0] = 14;
		pixel_array_in[3][1] = 60;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[25, 12, 23, 12],\n[46, 34, 48, 42],\n[25, 56, 5, 48],\n[6, 49, 1, 39]]");
		$display("Expect: 147, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 14;
		pixel_array_in[0][1] = 35;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 12;
		pixel_array_in[1][1] = 56;
		pixel_array_in[1][2] = 21;
		pixel_array_in[1][3] = 7;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 38;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 49;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 19;
		pixel_array_in[3][3] = 61;
		#10;
		
		$display("Input: \n[[3, 59, 36, 59],\n[36, 49, 33, 30],\n[47, 56, 55, 34],\n[37, 44, 2, 43]]");
		$display("Expect: 205, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 39;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 17;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 31;
		pixel_array_in[1][2] = 42;
		pixel_array_in[1][3] = 20;
		pixel_array_in[2][0] = 37;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 15;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 39;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 32;
		#10;
		
		$display("Input: \n[[56, 58, 12, 53],\n[28, 35, 42, 58],\n[10, 4, 20, 38],\n[13, 27, 1, 23]]");
		$display("Expect: 97, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 40;
		pixel_array_in[0][1] = 16;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 16;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 28;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 24;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 17;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[12, 20, 30, 2],\n[18, 58, 41, 48],\n[49, 42, 15, 2],\n[14, 60, 56, 52]]");
		$display("Expect: 158, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 43;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 26;
		pixel_array_in[0][3] = 34;
		pixel_array_in[1][0] = 23;
		pixel_array_in[1][1] = 42;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 34;
		pixel_array_in[2][0] = 9;
		pixel_array_in[2][1] = 25;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 59;
		pixel_array_in[3][1] = 54;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[14, 35, 30, 8],\n[12, 56, 21, 7],\n[15, 13, 38, 49],\n[49, 14, 19, 61]]");
		$display("Expect: 138, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 38;
		pixel_array_in[0][1] = 41;
		pixel_array_in[0][2] = 49;
		pixel_array_in[0][3] = 38;
		pixel_array_in[1][0] = 49;
		pixel_array_in[1][1] = 19;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 26;
		pixel_array_in[2][2] = 39;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 48;
		pixel_array_in[3][1] = 21;
		pixel_array_in[3][2] = 13;
		pixel_array_in[3][3] = 17;
		#10;
		
		$display("Input: \n[[39, 25, 7, 17],\n[47, 31, 42, 20],\n[37, 7, 0, 15],\n[41, 39, 15, 32]]");
		$display("Expect: 74, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 46;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 45;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 16;
		pixel_array_in[1][3] = 49;
		pixel_array_in[2][0] = 41;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 41;
		pixel_array_in[2][3] = 8;
		pixel_array_in[3][0] = 4;
		pixel_array_in[3][1] = 20;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 34;
		#10;
		
		$display("Input: \n[[40, 16, 48, 39],\n[57, 16, 22, 28],\n[42, 24, 23, 17],\n[52, 18, 3, 33]]");
		$display("Expect: 77, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 33;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 11;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 16;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 60;
		pixel_array_in[2][2] = 18;
		pixel_array_in[2][3] = 54;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 8;
		pixel_array_in[3][2] = 57;
		pixel_array_in[3][3] = 41;
		#10;
		
		$display("Input: \n[[43, 26, 26, 34],\n[23, 42, 56, 34],\n[9, 25, 19, 42],\n[59, 54, 6, 16]]");
		$display("Expect: 151, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 44;
		pixel_array_in[0][1] = 50;
		pixel_array_in[0][2] = 16;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 8;
		pixel_array_in[1][1] = 30;
		pixel_array_in[1][2] = 20;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 59;
		pixel_array_in[3][0] = 4;
		pixel_array_in[3][1] = 62;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[38, 41, 49, 38],\n[49, 19, 15, 6],\n[40, 26, 39, 18],\n[48, 21, 13, 17]]");
		$display("Expect: 94, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 28;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 38;
		pixel_array_in[0][3] = 23;
		pixel_array_in[1][0] = 41;
		pixel_array_in[1][1] = 31;
		pixel_array_in[1][2] = 42;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 62;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 56;
		pixel_array_in[2][3] = 29;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[15, 46, 21, 40],\n[45, 23, 16, 49],\n[41, 1, 41, 8],\n[4, 20, 7, 34]]");
		$display("Expect: 70, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 13;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 61;
		pixel_array_in[1][0] = 60;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 27;
		pixel_array_in[1][3] = 60;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 50;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[33, 17, 11, 45],\n[61, 12, 11, 16],\n[10, 60, 18, 54],\n[41, 8, 57, 41]]");
		$display("Expect: 97, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 58;
		pixel_array_in[0][1] = 34;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 38;
		pixel_array_in[1][2] = 47;
		pixel_array_in[1][3] = 42;
		pixel_array_in[2][0] = 27;
		pixel_array_in[2][1] = 31;
		pixel_array_in[2][2] = 24;
		pixel_array_in[2][3] = 27;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 15;
		pixel_array_in[3][2] = 5;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[44, 50, 16, 8],\n[8, 30, 20, 35],\n[31, 57, 23, 59],\n[4, 62, 36, 12]]");
		$display("Expect: 123, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 10;
		pixel_array_in[0][1] = 61;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 35;
		pixel_array_in[1][0] = 24;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 6;
		pixel_array_in[1][3] = 33;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[28, 40, 38, 23],\n[41, 31, 42, 6],\n[62, 36, 56, 29],\n[5, 44, 0, 20]]");
		$display("Expect: 173, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 29;
		pixel_array_in[0][3] = 50;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 20;
		pixel_array_in[1][3] = 28;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 19;
		pixel_array_in[2][2] = 60;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 35;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 57;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[53, 13, 19, 61],\n[60, 25, 27, 60],\n[24, 11, 44, 30],\n[50, 6, 42, 58]]");
		$display("Expect: 103, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 29;
		pixel_array_in[0][2] = 9;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 35;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 2;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 58;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 24;
		pixel_array_in[2][3] = 6;
		pixel_array_in[3][0] = 39;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 20;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[58, 34, 13, 41],\n[61, 38, 47, 42],\n[27, 31, 24, 27],\n[52, 15, 5, 12]]");
		$display("Expect: 148, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 20;
		pixel_array_in[0][2] = 2;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 14;
		pixel_array_in[1][1] = 15;
		pixel_array_in[1][2] = 12;
		pixel_array_in[1][3] = 37;
		pixel_array_in[2][0] = 26;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 27;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 29;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[10, 61, 14, 35],\n[24, 23, 6, 33],\n[14, 12, 42, 18],\n[17, 42, 7, 42]]");
		$display("Expect: 76, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 17;
		pixel_array_in[0][1] = 60;
		pixel_array_in[0][2] = 44;
		pixel_array_in[0][3] = 23;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 10;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 22;
		pixel_array_in[2][0] = 33;
		pixel_array_in[2][1] = 26;
		pixel_array_in[2][2] = 58;
		pixel_array_in[2][3] = 20;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 27;
		pixel_array_in[3][2] = 13;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[32, 32, 29, 50],\n[46, 60, 20, 28],\n[15, 19, 60, 1],\n[35, 58, 57, 12]]");
		$display("Expect: 165, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 20;
		pixel_array_in[0][1] = 44;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 28;
		pixel_array_in[1][0] = 8;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 42;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 18;
		pixel_array_in[2][3] = 8;
		pixel_array_in[3][0] = 26;
		pixel_array_in[3][1] = 19;
		pixel_array_in[3][2] = 25;
		pixel_array_in[3][3] = 9;
		#10;
		
		$display("Input: \n[[0, 29, 9, 8],\n[35, 49, 2, 48],\n[58, 23, 24, 6],\n[39, 48, 20, 7]]");
		$display("Expect: 89, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 14;
		pixel_array_in[0][1] = 4;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 62;
		pixel_array_in[1][2] = 46;
		pixel_array_in[1][3] = 37;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 34;
		pixel_array_in[3][0] = 47;
		pixel_array_in[3][1] = 17;
		pixel_array_in[3][2] = 1;
		pixel_array_in[3][3] = 25;
		#10;
		
		$display("Input: \n[[61, 20, 2, 15],\n[14, 15, 12, 37],\n[26, 40, 52, 27],\n[29, 29, 32, 27]]");
		$display("Expect: 126, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 11;
		pixel_array_in[0][2] = 58;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 23;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 41;
		pixel_array_in[2][0] = 16;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 20;
		pixel_array_in[3][0] = 60;
		pixel_array_in[3][1] = 61;
		pixel_array_in[3][2] = 38;
		pixel_array_in[3][3] = 26;
		#10;
		
		$display("Input: \n[[17, 60, 44, 23],\n[32, 10, 5, 22],\n[33, 26, 58, 20],\n[41, 27, 13, 33]]");
		$display("Expect: 91, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 36;
		pixel_array_in[0][2] = 36;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 8;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 18;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 34;
		pixel_array_in[2][2] = 25;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[20, 44, 4, 28],\n[8, 52, 56, 42],\n[31, 44, 18, 8],\n[26, 19, 25, 9]]");
		$display("Expect: 191, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 61;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 38;
		pixel_array_in[1][2] = 42;
		pixel_array_in[1][3] = 26;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 16;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 60;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[14, 4, 12, 2],\n[46, 62, 46, 37],\n[31, 40, 19, 34],\n[47, 17, 1, 25]]");
		$display("Expect: 187, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 37;
		pixel_array_in[0][2] = 42;
		pixel_array_in[0][3] = 22;
		pixel_array_in[1][0] = 27;
		pixel_array_in[1][1] = 55;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 49;
		pixel_array_in[2][1] = 31;
		pixel_array_in[2][2] = 16;
		pixel_array_in[2][3] = 13;
		pixel_array_in[3][0] = 14;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 15;
		#10;
		
		$display("Input: \n[[22, 11, 58, 44],\n[23, 49, 5, 41],\n[16, 7, 44, 20],\n[60, 61, 38, 26]]");
		$display("Expect: 97, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 50;
		pixel_array_in[0][1] = 38;
		pixel_array_in[0][2] = 29;
		pixel_array_in[0][3] = 16;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 31;
		pixel_array_in[1][3] = 58;
		pixel_array_in[2][0] = 52;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 13;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 11;
		pixel_array_in[3][1] = 10;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 19;
		#10;
		
		$display("Input: \n[[22, 36, 36, 53],\n[8, 12, 18, 44],\n[11, 34, 25, 25],\n[38, 45, 2, 20]]");
		$display("Expect: 85, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 60;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 54;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 18;
		pixel_array_in[1][2] = 41;
		pixel_array_in[1][3] = 11;
		pixel_array_in[2][0] = 35;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 48;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 34;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[29, 61, 7, 53],\n[44, 38, 42, 26],\n[15, 16, 5, 60],\n[25, 14, 48, 42]]");
		$display("Expect: 91, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 36;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 59;
		pixel_array_in[1][1] = 34;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 21;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 51;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 51;
		pixel_array_in[3][0] = 59;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 18;
		#10;
		
		$display("Input: \n[[21, 37, 42, 22],\n[27, 55, 36, 18],\n[49, 31, 16, 13],\n[14, 45, 56, 15]]");
		$display("Expect: 135, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 31;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 17;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 45;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 3;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 20;
		pixel_array_in[2][3] = 51;
		pixel_array_in[3][0] = 26;
		pixel_array_in[3][1] = 53;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 38;
		#10;
		
		$display("Input: \n[[50, 38, 29, 16],\n[22, 37, 31, 58],\n[52, 38, 13, 62],\n[11, 10, 3, 19]]");
		$display("Expect: 113, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 24;
		pixel_array_in[0][1] = 59;
		pixel_array_in[0][2] = 29;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 56;
		pixel_array_in[1][1] = 41;
		pixel_array_in[1][2] = 4;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 21;
		pixel_array_in[2][1] = 47;
		pixel_array_in[2][2] = 56;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 54;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[60, 26, 54, 18],\n[28, 18, 41, 11],\n[35, 3, 48, 55],\n[34, 6, 32, 58]]");
		$display("Expect: 107, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 11;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 6;
		pixel_array_in[0][3] = 27;
		pixel_array_in[1][0] = 56;
		pixel_array_in[1][1] = 34;
		pixel_array_in[1][2] = 52;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 44;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 15;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 47;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[36, 25, 34, 8],\n[59, 34, 25, 21],\n[0, 51, 7, 51],\n[59, 45, 32, 18]]");
		$display("Expect: 112, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 37;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 12;
		pixel_array_in[1][1] = 5;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 33;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 25;
		pixel_array_in[2][3] = 45;
		pixel_array_in[3][0] = 48;
		pixel_array_in[3][1] = 9;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 41;
		#10;
		
		$display("Input: \n[[31, 7, 7, 53],\n[17, 60, 45, 0],\n[3, 44, 20, 51],\n[26, 53, 17, 38]]");
		$display("Expect: 194, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 7;
		pixel_array_in[0][1] = 53;
		pixel_array_in[0][2] = 36;
		pixel_array_in[0][3] = 7;
		pixel_array_in[1][0] = 26;
		pixel_array_in[1][1] = 43;
		pixel_array_in[1][2] = 2;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 61;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 7;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 10;
		pixel_array_in[3][2] = 9;
		pixel_array_in[3][3] = 47;
		#10;
		
		$display("Input: \n[[24, 59, 29, 19],\n[56, 41, 4, 56],\n[21, 47, 56, 18],\n[15, 28, 54, 44]]");
		$display("Expect: 143, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 31;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 43;
		pixel_array_in[2][0] = 32;
		pixel_array_in[2][1] = 51;
		pixel_array_in[2][2] = 28;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 53;
		pixel_array_in[3][1] = 16;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[11, 48, 6, 27],\n[56, 34, 52, 17],\n[44, 44, 15, 62],\n[10, 47, 48, 20]]");
		$display("Expect: 138, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 38;
		pixel_array_in[0][1] = 49;
		pixel_array_in[0][2] = 5;
		pixel_array_in[0][3] = 31;
		pixel_array_in[1][0] = 30;
		pixel_array_in[1][1] = 34;
		pixel_array_in[1][2] = 61;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 24;
		pixel_array_in[2][2] = 27;
		pixel_array_in[2][3] = 34;
		pixel_array_in[3][0] = 33;
		pixel_array_in[3][1] = 39;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[29, 37, 51, 45],\n[12, 5, 5, 33],\n[47, 13, 25, 45],\n[48, 9, 42, 41]]");
		$display("Expect: 24, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 41;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 8;
		pixel_array_in[1][1] = 5;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 40;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 21;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 26;
		pixel_array_in[3][3] = 18;
		#10;
		
		$display("Input: \n[[7, 53, 36, 7],\n[26, 43, 2, 32],\n[31, 61, 49, 7],\n[23, 10, 9, 47]]");
		$display("Expect: 168, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 6;
		pixel_array_in[0][1] = 13;
		pixel_array_in[0][2] = 5;
		pixel_array_in[0][3] = 21;
		pixel_array_in[1][0] = 6;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 5;
		pixel_array_in[2][2] = 15;
		pixel_array_in[2][3] = 38;
		pixel_array_in[3][0] = 28;
		pixel_array_in[3][1] = 53;
		pixel_array_in[3][2] = 21;
		pixel_array_in[3][3] = 23;
		#10;
		
		$display("Input: \n[[31, 32, 19, 42],\n[11, 27, 30, 43],\n[32, 51, 28, 62],\n[53, 16, 15, 52]]");
		$display("Expect: 142, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 38;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 43;
		pixel_array_in[1][2] = 57;
		pixel_array_in[1][3] = 42;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 18;
		pixel_array_in[2][2] = 9;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 35;
		pixel_array_in[3][1] = 12;
		pixel_array_in[3][2] = 8;
		pixel_array_in[3][3] = 48;
		#10;
		
		$display("Input: \n[[38, 49, 5, 31],\n[30, 34, 61, 39],\n[43, 24, 27, 34],\n[33, 39, 2, 20]]");
		$display("Expect: 152, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 38;
		pixel_array_in[0][1] = 4;
		pixel_array_in[0][2] = 56;
		pixel_array_in[0][3] = 48;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 38;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 20;
		pixel_array_in[2][0] = 8;
		pixel_array_in[2][1] = 2;
		pixel_array_in[2][2] = 45;
		pixel_array_in[2][3] = 58;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 19;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 3;
		#10;
		
		$display("Input: \n[[57, 19, 41, 40],\n[8, 5, 25, 40],\n[22, 21, 43, 53],\n[32, 55, 26, 18]]");
		$display("Expect: 84, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 23;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 32;
		pixel_array_in[1][0] = 21;
		pixel_array_in[1][1] = 47;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 14;
		pixel_array_in[2][0] = 51;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 24;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 13;
		#10;
		
		$display("Input: \n[[6, 13, 5, 21],\n[6, 1, 15, 44],\n[11, 5, 15, 38],\n[28, 53, 21, 23]]");
		$display("Expect: 19, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 4;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 26;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 13;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 48;
		pixel_array_in[2][2] = 15;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 51;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 5;
		pixel_array_in[3][3] = 49;
		#10;
		
		$display("Input: \n[[38, 54, 12, 39],\n[32, 43, 57, 42],\n[43, 18, 9, 43],\n[35, 12, 8, 48]]");
		$display("Expect: 128, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 31;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 26;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 12;
		pixel_array_in[1][1] = 46;
		pixel_array_in[1][2] = 55;
		pixel_array_in[1][3] = 52;
		pixel_array_in[2][0] = 17;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 15;
		pixel_array_in[3][0] = 30;
		pixel_array_in[3][1] = 40;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 26;
		#10;
		
		$display("Input: \n[[38, 4, 56, 48],\n[9, 38, 37, 20],\n[8, 2, 45, 58],\n[41, 19, 15, 3]]");
		$display("Expect: 129, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 40;
		pixel_array_in[0][1] = 44;
		pixel_array_in[0][2] = 10;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 56;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 60;
		pixel_array_in[2][0] = 61;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 4;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 9;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 1;
		pixel_array_in[3][3] = 57;
		#10;
		
		$display("Input: \n[[22, 23, 51, 32],\n[21, 47, 0, 14],\n[51, 1, 24, 53],\n[41, 18, 27, 13]]");
		$display("Expect: 56, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 30;
		pixel_array_in[0][1] = 60;
		pixel_array_in[0][2] = 41;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 6;
		pixel_array_in[1][1] = 53;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 38;
		pixel_array_in[2][3] = 37;
		pixel_array_in[3][0] = 44;
		pixel_array_in[3][1] = 62;
		pixel_array_in[3][2] = 35;
		pixel_array_in[3][3] = 4;
		#10;
		
		$display("Input: \n[[4, 48, 7, 1],\n[28, 26, 36, 13],\n[57, 48, 15, 42],\n[51, 38, 5, 49]]");
		$display("Expect: 126, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 16;
		pixel_array_in[0][1] = 44;
		pixel_array_in[0][2] = 58;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 39;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 15;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 40;
		#10;
		
		$display("Input: \n[[31, 17, 26, 15],\n[12, 46, 55, 52],\n[17, 7, 47, 15],\n[30, 40, 36, 26]]");
		$display("Expect: 167, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 62;
		pixel_array_in[0][1] = 60;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 56;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 58;
		pixel_array_in[2][0] = 44;
		pixel_array_in[2][1] = 31;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 10;
		#10;
		
		$display("Input: \n[[40, 44, 10, 12],\n[56, 37, 3, 60],\n[61, 13, 4, 10],\n[9, 38, 1, 57]]");
		$display("Expect: 34, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 43;
		pixel_array_in[0][1] = 38;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 30;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 53;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 53;
		pixel_array_in[2][1] = 14;
		pixel_array_in[2][2] = 59;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 22;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 52;
		pixel_array_in[3][3] = 25;
		#10;
		
		$display("Input: \n[[30, 60, 41, 58],\n[6, 53, 56, 6],\n[39, 36, 38, 37],\n[44, 62, 35, 4]]");
		$display("Expect: 193, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 51;
		pixel_array_in[0][1] = 35;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 26;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 29;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 3;
		pixel_array_in[2][0] = 41;
		pixel_array_in[2][1] = 9;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 57;
		pixel_array_in[3][0] = 39;
		pixel_array_in[3][1] = 17;
		pixel_array_in[3][2] = 13;
		pixel_array_in[3][3] = 18;
		#10;
		
		$display("Input: \n[[16, 44, 58, 39],\n[39, 28, 39, 25],\n[12, 15, 47, 55],\n[25, 48, 11, 40]]");
		$display("Expect: 124, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 36;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 40;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 40;
		pixel_array_in[1][3] = 36;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 27;
		pixel_array_in[2][2] = 48;
		pixel_array_in[2][3] = 33;
		pixel_array_in[3][0] = 20;
		pixel_array_in[3][1] = 39;
		pixel_array_in[3][2] = 21;
		pixel_array_in[3][3] = 36;
		#10;
		
		$display("Input: \n[[62, 60, 13, 36],\n[61, 56, 5, 58],\n[44, 31, 0, 18],\n[19, 50, 59, 10]]");
		$display("Expect: 67, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 27;
		pixel_array_in[0][1] = 36;
		pixel_array_in[0][2] = 39;
		pixel_array_in[0][3] = 49;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 29;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 27;
		pixel_array_in[2][2] = 36;
		pixel_array_in[2][3] = 26;
		pixel_array_in[3][0] = 33;
		pixel_array_in[3][1] = 23;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[43, 38, 51, 30],\n[22, 53, 36, 17],\n[53, 14, 59, 1],\n[22, 18, 52, 25]]");
		$display("Expect: 171, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 9;
		pixel_array_in[0][2] = 62;
		pixel_array_in[0][3] = 13;
		pixel_array_in[1][0] = 36;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 1;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 41;
		pixel_array_in[2][1] = 20;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 55;
		#10;
		
		$display("Input: \n[[51, 35, 23, 26],\n[46, 29, 11, 3],\n[41, 9, 54, 57],\n[39, 17, 13, 18]]");
		$display("Expect: 99, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 5;
		pixel_array_in[0][1] = 22;
		pixel_array_in[0][2] = 1;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 30;
		pixel_array_in[1][2] = 41;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 35;
		pixel_array_in[2][1] = 19;
		pixel_array_in[2][2] = 40;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 50;
		pixel_array_in[3][1] = 62;
		pixel_array_in[3][2] = 8;
		pixel_array_in[3][3] = 61;
		#10;
		
		$display("Input: \n[[32, 17, 36, 15],\n[40, 60, 40, 36],\n[57, 27, 48, 33],\n[20, 39, 21, 36]]");
		$display("Expect: 183, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 54;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 53;
		pixel_array_in[1][1] = 46;
		pixel_array_in[1][2] = 28;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 49;
		pixel_array_in[2][1] = 25;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 48;
		pixel_array_in[3][0] = 51;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 8;
		#10;
		
		$display("Input: \n[[27, 36, 39, 49],\n[57, 29, 13, 25],\n[22, 27, 36, 26],\n[33, 23, 3, 6]]");
		$display("Expect: 102, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 20;
		pixel_array_in[0][2] = 35;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 51;
		pixel_array_in[1][1] = 3;
		pixel_array_in[1][2] = 61;
		pixel_array_in[1][3] = 2;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 39;
		pixel_array_in[2][2] = 37;
		pixel_array_in[2][3] = 33;
		pixel_array_in[3][0] = 35;
		pixel_array_in[3][1] = 2;
		pixel_array_in[3][2] = 35;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[29, 9, 62, 13],\n[36, 45, 1, 44],\n[41, 20, 5, 42],\n[19, 26, 17, 55]]");
		$display("Expect: 52, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 51;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 28;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 6;
		pixel_array_in[1][2] = 6;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 46;
		pixel_array_in[2][3] = 45;
		pixel_array_in[3][0] = 33;
		pixel_array_in[3][1] = 35;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[5, 22, 1, 18],\n[0, 30, 41, 44],\n[35, 19, 40, 44],\n[50, 62, 8, 61]]");
		$display("Expect: 136, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 55;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 51;
		pixel_array_in[1][0] = 33;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 4;
		pixel_array_in[2][3] = 29;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 9;
		#10;
		
		$display("Input: \n[[54, 32, 12, 0],\n[53, 46, 28, 39],\n[49, 25, 43, 48],\n[51, 34, 51, 8]]");
		$display("Expect: 136, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 16;
		pixel_array_in[0][3] = 47;
		pixel_array_in[1][0] = 36;
		pixel_array_in[1][1] = 51;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 30;
		pixel_array_in[2][0] = 7;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 55;
		pixel_array_in[2][3] = 52;
		pixel_array_in[3][0] = 39;
		pixel_array_in[3][1] = 20;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 46;
		#10;
		
		$display("Input: \n[[0, 20, 35, 59],\n[51, 3, 61, 2],\n[43, 39, 37, 33],\n[35, 2, 35, 60]]");
		$display("Expect: 148, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 35;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 7;
		pixel_array_in[1][1] = 57;
		pixel_array_in[1][2] = 45;
		pixel_array_in[1][3] = 41;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 12;
		pixel_array_in[2][3] = 59;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[51, 10, 51, 28],\n[10, 6, 6, 29],\n[30, 40, 46, 45],\n[33, 35, 55, 58]]");
		$display("Expect: 89, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 59;
		pixel_array_in[0][1] = 59;
		pixel_array_in[0][2] = 29;
		pixel_array_in[0][3] = 3;
		pixel_array_in[1][0] = 39;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 8;
		pixel_array_in[2][1] = 31;
		pixel_array_in[2][2] = 32;
		pixel_array_in[2][3] = 45;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 23;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[21, 55, 21, 51],\n[33, 0, 33, 25],\n[42, 7, 4, 29],\n[52, 6, 55, 9]]");
		$display("Expect: 20, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 3;
		pixel_array_in[0][1] = 22;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 29;
		pixel_array_in[1][0] = 15;
		pixel_array_in[1][1] = 41;
		pixel_array_in[1][2] = 40;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 26;
		pixel_array_in[2][1] = 8;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 21;
		pixel_array_in[3][1] = 21;
		pixel_array_in[3][2] = 30;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[19, 17, 16, 47],\n[36, 51, 22, 30],\n[7, 45, 55, 52],\n[39, 20, 32, 46]]");
		$display("Expect: 191, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 54;
		pixel_array_in[1][0] = 51;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 46;
		pixel_array_in[1][3] = 41;
		pixel_array_in[2][0] = 9;
		pixel_array_in[2][1] = 5;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 58;
		pixel_array_in[3][0] = 33;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 54;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[29, 25, 35, 12],\n[7, 57, 45, 41],\n[0, 44, 12, 59],\n[31, 6, 17, 60]]");
		$display("Expect: 175, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 20;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 52;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 34;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 62;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 12;
		pixel_array_in[3][0] = 6;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[59, 59, 29, 3],\n[39, 12, 0, 47],\n[8, 31, 32, 45],\n[42, 42, 23, 7]]");
		$display("Expect: 55, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 36;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 56;
		pixel_array_in[1][1] = 2;
		pixel_array_in[1][2] = 27;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 51;
		pixel_array_in[2][1] = 33;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 22;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 24;
		#10;
		
		$display("Input: \n[[3, 22, 19, 29],\n[15, 41, 40, 46],\n[26, 8, 57, 3],\n[21, 21, 30, 27]]");
		$display("Expect: 160, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 34;
		pixel_array_in[0][1] = 60;
		pixel_array_in[0][2] = 31;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 48;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 52;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 16;
		pixel_array_in[2][2] = 13;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 9;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[8, 26, 52, 54],\n[51, 45, 46, 41],\n[9, 5, 44, 58],\n[33, 25, 54, 44]]");
		$display("Expect: 134, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 38;
		pixel_array_in[0][3] = 51;
		pixel_array_in[1][0] = 49;
		pixel_array_in[1][1] = 62;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 34;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 40;
		pixel_array_in[2][3] = 27;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 46;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 28;
		#10;
		
		$display("Input: \n[[20, 45, 30, 44],\n[52, 32, 34, 29],\n[1, 62, 47, 12],\n[6, 44, 12, 39]]");
		$display("Expect: 191, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 18;
		pixel_array_in[0][1] = 9;
		pixel_array_in[0][2] = 39;
		pixel_array_in[0][3] = 56;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 8;
		pixel_array_in[1][3] = 54;
		pixel_array_in[2][0] = 54;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 29;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 46;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[36, 45, 23, 25],\n[56, 2, 27, 39],\n[51, 33, 49, 22],\n[17, 59, 45, 24]]");
		$display("Expect: 94, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 16;
		pixel_array_in[0][2] = 9;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 23;
		pixel_array_in[1][1] = 20;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 21;
		pixel_array_in[2][0] = 34;
		pixel_array_in[2][1] = 8;
		pixel_array_in[2][2] = 12;
		pixel_array_in[2][3] = 52;
		pixel_array_in[3][0] = 50;
		pixel_array_in[3][1] = 47;
		pixel_array_in[3][2] = 10;
		pixel_array_in[3][3] = 13;
		#10;
		
		$display("Input: \n[[34, 60, 31, 2],\n[47, 48, 39, 52],\n[31, 16, 13, 10],\n[15, 45, 9, 35]]");
		$display("Expect: 108, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 5;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 57;
		pixel_array_in[1][2] = 55;
		pixel_array_in[1][3] = 10;
		pixel_array_in[2][0] = 33;
		pixel_array_in[2][1] = 48;
		pixel_array_in[2][2] = 28;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 52;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[29, 18, 38, 51],\n[49, 62, 37, 34],\n[40, 32, 40, 27],\n[46, 46, 7, 28]]");
		$display("Expect: 182, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[18, 9, 39, 56],\n[11, 28, 8, 54],\n[54, 45, 42, 29],\n[32, 50, 46, 6]]");
		$display("Expect: 116, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[1, 16, 9, 40],\n[23, 20, 22, 21],\n[34, 8, 12, 52],\n[50, 47, 10, 13]]");
		$display("Expect: 50, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[5, 58, 52, 42],\n[31, 57, 55, 10],\n[33, 48, 28, 1],\n[15, 52, 61, 1]]");
		$display("Expect: 197, Result: %d", pixel_out);
		$display("");
		#10;
		
		
		$display("Finishing Sim"); //print nice message
		$finish;
		
    end
endmodule //counter_tb

`default_nettype wire