`timescale 1ns / 1ps
`default_nettype none

module kernel_3_tb;

    //make logics for inputs and outputs!
    logic clk_in;
    logic rst_in;
    logic valid_in;
    logic [5:0] pixel_array_in [3:0][3:0];
    logic [8:0] pixel_out;

    kernel_3 uut (
        .clk_in(clk_in),
        .p(pixel_array_in),
        .pixel_out(pixel_out)
    );
    always begin
        #5;  //every 5 ns switch...so period of clock is 10 ns...100 MHz clock
        clk_in = !clk_in;
    end

    //initial block...this is our test simulation
    initial begin

		$dumpfile("test/kernel_3.vcd"); //file to store value change dump (vcd)
		$dumpvars(0,kernel_3_tb); //store everything at the current level and below
		$display("Starting Sim"); //print nice message
		clk_in = 0; //initialize clk (super important)
		rst_in = 0; //initialize rst (super important)
		
		#10;  //wait a little bit of time at beginning
		rst_in = 1; //reset system
		#10; //hold high for a few clock cycles
		rst_in=0;
		
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 0;
		#10;
		
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 32;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 32;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 32;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 32;
		#10;
		
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 63;
		#10;
		
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 63;
		#10;
		
		$display("Input: \n[[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0]]");
		$display("Expect: 0, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Input: \n[[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32]]");
		$display("Expect: 128, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 5;
		pixel_array_in[0][2] = 60;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 2;
		pixel_array_in[1][2] = 59;
		pixel_array_in[1][3] = 54;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 43;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 11;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63]]");
		$display("Expect: 252, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 12;
		pixel_array_in[0][1] = 36;
		pixel_array_in[0][2] = 33;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 42;
		pixel_array_in[1][1] = 13;
		pixel_array_in[1][2] = 34;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 35;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 38;
		pixel_array_in[3][0] = 30;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 61;
		#10;
		
		$display("Input: \n[[63, 0, 0, 63],\n[0, 63, 63, 0],\n[0, 63, 63, 0],\n[63, 0, 0, 63]]");
		$display("Expect: 384>val>255, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 11;
		pixel_array_in[0][2] = 28;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 18;
		pixel_array_in[1][1] = 42;
		pixel_array_in[1][2] = 48;
		pixel_array_in[1][3] = 55;
		pixel_array_in[2][0] = 7;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 26;
		pixel_array_in[2][3] = 37;
		pixel_array_in[3][0] = 1;
		pixel_array_in[3][1] = 29;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[0, 63, 63, 0],\n[63, 0, 0, 63],\n[63, 0, 0, 63],\n[0, 63, 63, 0]]");
		$display("Expect: val>383, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 20;
		pixel_array_in[0][1] = 1;
		pixel_array_in[0][2] = 60;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 21;
		pixel_array_in[1][3] = 55;
		pixel_array_in[2][0] = 49;
		pixel_array_in[2][1] = 18;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 20;
		pixel_array_in[3][3] = 9;
		#10;
		
		$display("Input: \n[[32, 5, 60, 18],\n[57, 2, 59, 54],\n[31, 43, 30, 1],\n[15, 11, 36, 39]]");
		$display("Expect: 66, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 30;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 35;
		pixel_array_in[1][0] = 54;
		pixel_array_in[1][1] = 2;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 3;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 30;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 5;
		pixel_array_in[3][2] = 18;
		pixel_array_in[3][3] = 37;
		#10;
		
		$display("Input: \n[[12, 36, 33, 10],\n[42, 13, 34, 56],\n[35, 45, 61, 38],\n[30, 55, 45, 61]]");
		$display("Expect: 80, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 30;
		pixel_array_in[0][1] = 39;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 54;
		pixel_array_in[1][1] = 9;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 51;
		pixel_array_in[2][0] = 9;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 11;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 20;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 62;
		pixel_array_in[3][3] = 5;
		#10;
		
		$display("Input: \n[[22, 11, 28, 40],\n[18, 42, 48, 55],\n[7, 44, 26, 37],\n[1, 29, 56, 60]]");
		$display("Expect: 186, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 47;
		pixel_array_in[0][1] = 5;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 2;
		pixel_array_in[1][2] = 14;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 53;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 2;
		pixel_array_in[3][0] = 51;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 51;
		#10;
		
		$display("Input: \n[[20, 1, 60, 19],\n[11, 35, 21, 55],\n[49, 18, 30, 53],\n[25, 32, 20, 9]]");
		$display("Expect: 124, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 34;
		pixel_array_in[0][1] = 27;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 51;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 62;
		pixel_array_in[1][2] = 34;
		pixel_array_in[1][3] = 13;
		pixel_array_in[2][0] = 33;
		pixel_array_in[2][1] = 20;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 29;
		pixel_array_in[3][0] = 28;
		pixel_array_in[3][1] = 61;
		pixel_array_in[3][2] = 46;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[30, 52, 52, 35],\n[54, 2, 3, 3],\n[39, 30, 42, 49],\n[25, 5, 18, 37]]");
		$display("Expect: 7, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 60;
		pixel_array_in[0][1] = 6;
		pixel_array_in[0][2] = 31;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 8;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 2;
		pixel_array_in[2][2] = 35;
		pixel_array_in[2][3] = 28;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 47;
		pixel_array_in[3][3] = 30;
		#10;
		
		$display("Input: \n[[30, 39, 51, 39],\n[54, 9, 10, 51],\n[9, 12, 11, 3],\n[20, 50, 62, 5]]");
		$display("Expect: 11, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 50;
		pixel_array_in[0][1] = 50;
		pixel_array_in[0][2] = 62;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 21;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 49;
		pixel_array_in[1][3] = 57;
		pixel_array_in[2][0] = 51;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 6;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 6;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 31;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[47, 5, 23, 59],\n[10, 2, 14, 4],\n[53, 10, 17, 2],\n[51, 45, 42, 51]]");
		$display("Expect: 16, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 39;
		pixel_array_in[0][2] = 22;
		pixel_array_in[0][3] = 35;
		pixel_array_in[1][0] = 1;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 19;
		pixel_array_in[2][1] = 53;
		pixel_array_in[2][2] = 21;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 3;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 5;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[34, 27, 19, 51],\n[13, 62, 34, 13],\n[33, 20, 54, 29],\n[28, 61, 46, 33]]");
		$display("Expect: 220, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 42;
		pixel_array_in[0][1] = 36;
		pixel_array_in[0][2] = 37;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 53;
		pixel_array_in[1][2] = 35;
		pixel_array_in[1][3] = 1;
		pixel_array_in[2][0] = 49;
		pixel_array_in[2][1] = 4;
		pixel_array_in[2][2] = 15;
		pixel_array_in[2][3] = 4;
		pixel_array_in[3][0] = 49;
		pixel_array_in[3][1] = 62;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[60, 6, 31, 42],\n[31, 1, 8, 38],\n[47, 2, 35, 28],\n[42, 28, 47, 30]]");
		$display("Expect: val>383, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 48;
		pixel_array_in[0][1] = 8;
		pixel_array_in[0][2] = 53;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 52;
		pixel_array_in[1][1] = 40;
		pixel_array_in[1][2] = 52;
		pixel_array_in[1][3] = 60;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 56;
		pixel_array_in[2][3] = 59;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 10;
		#10;
		
		$display("Input: \n[[50, 50, 62, 36],\n[21, 52, 49, 57],\n[51, 3, 6, 3],\n[6, 44, 31, 20]]");
		$display("Expect: 166, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 39;
		pixel_array_in[0][1] = 31;
		pixel_array_in[0][2] = 2;
		pixel_array_in[0][3] = 27;
		pixel_array_in[1][0] = 24;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 41;
		pixel_array_in[1][3] = 41;
		pixel_array_in[2][0] = 2;
		pixel_array_in[2][1] = 58;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 14;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[9, 39, 22, 35],\n[1, 52, 15, 4],\n[19, 53, 21, 41],\n[3, 38, 5, 42]]");
		$display("Expect: 197, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 35;
		pixel_array_in[0][1] = 41;
		pixel_array_in[0][2] = 25;
		pixel_array_in[0][3] = 14;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 53;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 34;
		pixel_array_in[2][0] = 28;
		pixel_array_in[2][1] = 46;
		pixel_array_in[2][2] = 46;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 45;
		#10;
		
		$display("Input: \n[[42, 36, 37, 53],\n[58, 53, 35, 1],\n[49, 4, 15, 4],\n[49, 62, 55, 33]]");
		$display("Expect: 159, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 31;
		pixel_array_in[0][1] = 60;
		pixel_array_in[0][2] = 41;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 11;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 58;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 34;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 47;
		pixel_array_in[3][1] = 60;
		pixel_array_in[3][2] = 25;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[48, 8, 53, 40],\n[52, 40, 52, 60],\n[57, 10, 56, 59],\n[13, 14, 45, 10]]");
		$display("Expect: 152, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 10;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 47;
		pixel_array_in[0][3] = 13;
		pixel_array_in[1][0] = 24;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 21;
		pixel_array_in[1][3] = 53;
		pixel_array_in[2][0] = 6;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 34;
		pixel_array_in[2][3] = 51;
		pixel_array_in[3][0] = 20;
		pixel_array_in[3][1] = 12;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Input: \n[[39, 31, 2, 27],\n[24, 0, 41, 41],\n[2, 58, 61, 41],\n[14, 32, 29, 16]]");
		$display("Expect: 70, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 60;
		pixel_array_in[0][1] = 36;
		pixel_array_in[0][2] = 26;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 45;
		pixel_array_in[2][1] = 54;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 37;
		pixel_array_in[3][1] = 9;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 61;
		#10;
		
		$display("Input: \n[[35, 41, 25, 14],\n[0, 53, 0, 34],\n[28, 46, 46, 55],\n[52, 55, 11, 45]]");
		$display("Expect: 184, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 26;
		pixel_array_in[0][1] = 2;
		pixel_array_in[0][2] = 8;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 33;
		pixel_array_in[1][1] = 40;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 30;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 41;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 36;
		#10;
		
		$display("Input: \n[[31, 60, 41, 15],\n[46, 11, 56, 39],\n[58, 13, 34, 39],\n[47, 60, 25, 56]]");
		$display("Expect: 54, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 27;
		pixel_array_in[0][1] = 11;
		pixel_array_in[0][2] = 54;
		pixel_array_in[0][3] = 14;
		pixel_array_in[1][0] = 54;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 8;
		pixel_array_in[1][3] = 31;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 1;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[10, 25, 47, 13],\n[24, 54, 21, 53],\n[6, 55, 34, 51],\n[20, 12, 45, 0]]");
		$display("Expect: 207, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 62;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 26;
		pixel_array_in[0][3] = 61;
		pixel_array_in[1][0] = 49;
		pixel_array_in[1][1] = 6;
		pixel_array_in[1][2] = 23;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 21;
		pixel_array_in[2][1] = 16;
		pixel_array_in[2][2] = 11;
		pixel_array_in[2][3] = 51;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 33;
		pixel_array_in[3][3] = 49;
		#10;
		
		$display("Input: \n[[60, 36, 26, 12],\n[46, 32, 50, 12],\n[45, 54, 42, 39],\n[37, 9, 61, 61]]");
		$display("Expect: 159, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 13;
		pixel_array_in[0][2] = 9;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 48;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 62;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 48;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 45;
		#10;
		
		$display("Input: \n[[26, 2, 8, 59],\n[33, 40, 37, 30],\n[60, 41, 44, 44],\n[40, 59, 51, 36]]");
		$display("Expect: 169, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 24;
		pixel_array_in[0][2] = 58;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 31;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 25;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 47;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 10;
		#10;
		
		$display("Input: \n[[27, 11, 54, 14],\n[54, 60, 8, 31],\n[5, 44, 1, 30],\n[5, 37, 15, 60]]");
		$display("Expect: 196, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 24;
		pixel_array_in[0][2] = 36;
		pixel_array_in[0][3] = 61;
		pixel_array_in[1][0] = 8;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 54;
		pixel_array_in[1][3] = 22;
		pixel_array_in[2][0] = 45;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 3;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 53;
		#10;
		
		$display("Input: \n[[62, 28, 26, 61],\n[49, 6, 23, 46],\n[21, 16, 11, 51],\n[13, 50, 33, 49]]");
		$display("Expect: 21, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 31;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 33;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 28;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 19;
		pixel_array_in[3][2] = 33;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[9, 13, 9, 36],\n[48, 25, 30, 32],\n[24, 62, 61, 48],\n[13, 48, 60, 45]]");
		$display("Expect: 134, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 44;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 37;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 26;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 35;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[57, 24, 58, 33],\n[58, 31, 25, 62],\n[57, 17, 25, 42],\n[47, 37, 2, 10]]");
		$display("Expect: 96, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 5;
		pixel_array_in[0][1] = 53;
		pixel_array_in[0][2] = 43;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 43;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 18;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 30;
		pixel_array_in[2][2] = 56;
		pixel_array_in[2][3] = 57;
		pixel_array_in[3][0] = 56;
		pixel_array_in[3][1] = 61;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 34;
		#10;
		
		$display("Input: \n[[61, 24, 36, 61],\n[8, 27, 54, 22],\n[45, 55, 7, 41],\n[46, 3, 7, 53]]");
		$display("Expect: 154, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 29;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 24;
		pixel_array_in[1][0] = 34;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 47;
		pixel_array_in[1][3] = 37;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 52;
		pixel_array_in[2][2] = 40;
		pixel_array_in[2][3] = 21;
		pixel_array_in[3][0] = 6;
		pixel_array_in[3][1] = 19;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[31, 18, 33, 41],\n[38, 33, 28, 18],\n[11, 7, 44, 1],\n[5, 19, 33, 7]]");
		$display("Expect: 116, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 6;
		pixel_array_in[0][1] = 41;
		pixel_array_in[0][2] = 27;
		pixel_array_in[0][3] = 62;
		pixel_array_in[1][0] = 53;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 59;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 20;
		pixel_array_in[2][3] = 12;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 43;
		pixel_array_in[3][2] = 30;
		pixel_array_in[3][3] = 19;
		#10;
		
		$display("Input: \n[[44, 54, 4, 37],\n[11, 50, 26, 44],\n[60, 40, 52, 44],\n[35, 50, 2, 33]]");
		$display("Expect: 185, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 50;
		pixel_array_in[0][1] = 30;
		pixel_array_in[0][2] = 33;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 55;
		pixel_array_in[1][1] = 3;
		pixel_array_in[1][2] = 48;
		pixel_array_in[1][3] = 3;
		pixel_array_in[2][0] = 53;
		pixel_array_in[2][1] = 24;
		pixel_array_in[2][2] = 53;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[5, 53, 43, 58],\n[43, 23, 18, 35],\n[22, 30, 56, 57],\n[56, 61, 12, 34]]");
		$display("Expect: 82, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 41;
		pixel_array_in[0][1] = 16;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 43;
		pixel_array_in[1][0] = 3;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 62;
		pixel_array_in[1][3] = 59;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 59;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 60;
		pixel_array_in[3][1] = 22;
		pixel_array_in[3][2] = 49;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[22, 29, 13, 24],\n[34, 27, 47, 37],\n[39, 52, 40, 21],\n[6, 19, 36, 52]]");
		$display("Expect: 143, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 46;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 43;
		pixel_array_in[0][3] = 22;
		pixel_array_in[1][0] = 14;
		pixel_array_in[1][1] = 9;
		pixel_array_in[1][2] = 52;
		pixel_array_in[1][3] = 10;
		pixel_array_in[2][0] = 3;
		pixel_array_in[2][1] = 5;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 17;
		pixel_array_in[3][2] = 26;
		pixel_array_in[3][3] = 25;
		#10;
		
		$display("Input: \n[[6, 41, 27, 62],\n[53, 25, 10, 59],\n[30, 36, 20, 12],\n[13, 43, 30, 19]]");
		$display("Expect: 80, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 8;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 46;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 13;
		pixel_array_in[2][1] = 19;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 16;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 62;
		#10;
		
		$display("Input: \n[[50, 30, 33, 58],\n[55, 3, 48, 3],\n[53, 24, 53, 30],\n[38, 55, 2, 58]]");
		$display("Expect: 46, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 11;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 7;
		pixel_array_in[1][3] = 10;
		pixel_array_in[2][0] = 37;
		pixel_array_in[2][1] = 19;
		pixel_array_in[2][2] = 58;
		pixel_array_in[2][3] = 19;
		pixel_array_in[3][0] = 48;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[41, 16, 0, 43],\n[3, 1, 62, 59],\n[30, 59, 42, 1],\n[60, 22, 49, 58]]");
		$display("Expect: 94, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 27;
		pixel_array_in[0][1] = 30;
		pixel_array_in[0][2] = 3;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 51;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 38;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 21;
		pixel_array_in[2][2] = 38;
		pixel_array_in[2][3] = 23;
		pixel_array_in[3][0] = 1;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[46, 48, 43, 22],\n[14, 9, 52, 10],\n[3, 5, 17, 25],\n[61, 17, 26, 25]]");
		$display("Expect: 55, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 14;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 6;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 27;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 28;
		pixel_array_in[3][3] = 54;
		#10;
		
		$display("Input: \n[[25, 8, 45, 12],\n[31, 28, 46, 12],\n[13, 19, 44, 3],\n[16, 45, 2, 62]]");
		$display("Expect: 127, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 47;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 15;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 9;
		pixel_array_in[1][3] = 54;
		pixel_array_in[2][0] = 53;
		pixel_array_in[2][1] = 60;
		pixel_array_in[2][2] = 36;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 26;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 28;
		#10;
		
		$display("Input: \n[[9, 28, 11, 8],\n[9, 50, 7, 10],\n[37, 19, 58, 19],\n[48, 37, 51, 56]]");
		$display("Expect: 165, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 7;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 56;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 39;
		pixel_array_in[1][2] = 51;
		pixel_array_in[1][3] = 5;
		pixel_array_in[2][0] = 8;
		pixel_array_in[2][1] = 24;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 50;
		pixel_array_in[3][0] = 62;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 23;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[27, 30, 3, 0],\n[51, 54, 38, 18],\n[15, 21, 38, 23],\n[1, 14, 48, 1]]");
		$display("Expect: 192, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 30;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 60;
		pixel_array_in[1][1] = 9;
		pixel_array_in[1][2] = 40;
		pixel_array_in[1][3] = 14;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 16;
		pixel_array_in[2][2] = 26;
		pixel_array_in[2][3] = 54;
		pixel_array_in[3][0] = 24;
		pixel_array_in[3][1] = 29;
		pixel_array_in[3][2] = 44;
		pixel_array_in[3][3] = 41;
		#10;
		
		$display("Input: \n[[1, 28, 21, 39],\n[14, 37, 6, 62],\n[27, 17, 47, 36],\n[10, 28, 28, 54]]");
		$display("Expect: 117, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 49;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 31;
		pixel_array_in[0][3] = 26;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 27;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 59;
		pixel_array_in[2][2] = 21;
		pixel_array_in[2][3] = 52;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 7;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 28;
		#10;
		
		$display("Input: \n[[47, 19, 15, 18],\n[31, 49, 9, 54],\n[53, 60, 36, 39],\n[26, 38, 11, 28]]");
		$display("Expect: 185, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 3;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 48;
		pixel_array_in[1][0] = 34;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 33;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 19;
		pixel_array_in[2][2] = 34;
		pixel_array_in[2][3] = 8;
		pixel_array_in[3][0] = 22;
		pixel_array_in[3][1] = 16;
		pixel_array_in[3][2] = 58;
		pixel_array_in[3][3] = 19;
		#10;
		
		$display("Input: \n[[7, 7, 56, 58],\n[10, 39, 51, 5],\n[8, 24, 47, 50],\n[62, 42, 23, 60]]");
		$display("Expect: 172, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 13;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 37;
		pixel_array_in[1][0] = 40;
		pixel_array_in[1][1] = 42;
		pixel_array_in[1][2] = 9;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 3;
		pixel_array_in[2][1] = 26;
		pixel_array_in[2][2] = 35;
		pixel_array_in[2][3] = 4;
		pixel_array_in[3][0] = 49;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 54;
		#10;
		
		$display("Input: \n[[53, 30, 19, 25],\n[60, 9, 40, 14],\n[11, 16, 26, 54],\n[24, 29, 44, 41]]");
		$display("Expect: 48, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 11;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 62;
		pixel_array_in[1][0] = 16;
		pixel_array_in[1][1] = 39;
		pixel_array_in[1][2] = 49;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 61;
		pixel_array_in[2][2] = 2;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 41;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[49, 0, 31, 26],\n[32, 1, 27, 38],\n[5, 59, 21, 52],\n[15, 7, 45, 28]]");
		$display("Expect: 60, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 38;
		pixel_array_in[0][1] = 53;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 15;
		pixel_array_in[1][1] = 20;
		pixel_array_in[1][2] = 55;
		pixel_array_in[1][3] = 45;
		pixel_array_in[2][0] = 33;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 58;
		pixel_array_in[2][3] = 6;
		pixel_array_in[3][0] = 9;
		pixel_array_in[3][1] = 11;
		pixel_array_in[3][2] = 19;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[29, 3, 55, 48],\n[34, 33, 37, 33],\n[5, 19, 34, 8],\n[22, 16, 58, 19]]");
		$display("Expect: 132, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 4;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 18;
		pixel_array_in[0][3] = 34;
		pixel_array_in[1][0] = 30;
		pixel_array_in[1][1] = 26;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 29;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 34;
		pixel_array_in[3][0] = 59;
		pixel_array_in[3][1] = 8;
		pixel_array_in[3][2] = 37;
		pixel_array_in[3][3] = 53;
		#10;
		
		$display("Input: \n[[13, 26, 48, 37],\n[40, 42, 9, 35],\n[3, 26, 35, 4],\n[49, 44, 61, 54]]");
		$display("Expect: 134, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 34;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 58;
		pixel_array_in[1][2] = 49;
		pixel_array_in[1][3] = 42;
		pixel_array_in[2][0] = 35;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 45;
		pixel_array_in[2][3] = 59;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 46;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 49;
		#10;
		
		$display("Input: \n[[11, 0, 55, 62],\n[16, 39, 49, 46],\n[22, 61, 2, 41],\n[5, 38, 41, 7]]");
		$display("Expect: 187, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 46;
		pixel_array_in[0][3] = 11;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 31;
		pixel_array_in[2][0] = 19;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 9;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 55;
		pixel_array_in[3][1] = 11;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[38, 53, 23, 55],\n[15, 20, 55, 45],\n[33, 44, 58, 6],\n[9, 11, 19, 58]]");
		$display("Expect: 126, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 47;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 7;
		pixel_array_in[1][1] = 48;
		pixel_array_in[1][2] = 52;
		pixel_array_in[1][3] = 8;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 28;
		pixel_array_in[2][2] = 8;
		pixel_array_in[2][3] = 60;
		pixel_array_in[3][0] = 30;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 28;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[4, 52, 18, 34],\n[30, 26, 22, 44],\n[22, 29, 7, 34],\n[59, 8, 37, 53]]");
		$display("Expect: 91, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 50;
		pixel_array_in[0][2] = 61;
		pixel_array_in[0][3] = 3;
		pixel_array_in[1][0] = 52;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 41;
		pixel_array_in[1][3] = 49;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 37;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 21;
		pixel_array_in[3][2] = 24;
		pixel_array_in[3][3] = 28;
		#10;
		
		$display("Input: \n[[0, 19, 13, 34],\n[22, 58, 49, 42],\n[35, 11, 45, 59],\n[42, 46, 29, 49]]");
		$display("Expect: 209, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 37;
		pixel_array_in[0][1] = 20;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 21;
		pixel_array_in[1][0] = 56;
		pixel_array_in[1][1] = 9;
		pixel_array_in[1][2] = 14;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 18;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 41;
		pixel_array_in[3][2] = 43;
		pixel_array_in[3][3] = 38;
		#10;
		
		$display("Input: \n[[0, 54, 46, 11],\n[58, 45, 39, 31],\n[19, 35, 9, 32],\n[55, 11, 56, 35]]");
		$display("Expect: 159, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 34;
		pixel_array_in[0][1] = 24;
		pixel_array_in[0][2] = 22;
		pixel_array_in[0][3] = 54;
		pixel_array_in[1][0] = 21;
		pixel_array_in[1][1] = 19;
		pixel_array_in[1][2] = 7;
		pixel_array_in[1][3] = 22;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 59;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[0, 47, 45, 8],\n[7, 48, 52, 8],\n[14, 28, 8, 60],\n[30, 45, 28, 42]]");
		$display("Expect: 186, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 5;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 61;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 41;
		pixel_array_in[1][2] = 54;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 45;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 7;
		pixel_array_in[3][1] = 62;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 25;
		#10;
		
		$display("Input: \n[[22, 50, 61, 3],\n[52, 33, 41, 49],\n[14, 32, 17, 37],\n[10, 21, 24, 28]]");
		$display("Expect: 124, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 25;
		pixel_array_in[1][1] = 29;
		pixel_array_in[1][2] = 62;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 14;
		pixel_array_in[2][2] = 51;
		pixel_array_in[2][3] = 54;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 48;
		#10;
		
		$display("Input: \n[[37, 20, 51, 21],\n[56, 9, 14, 18],\n[1, 18, 5, 25],\n[25, 41, 43, 38]]");
		$display("Expect: 26, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 5;
		pixel_array_in[0][2] = 17;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 37;
		pixel_array_in[1][1] = 44;
		pixel_array_in[1][2] = 44;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 23;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 15;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 54;
		#10;
		
		$display("Input: \n[[34, 24, 22, 54],\n[21, 19, 7, 22],\n[12, 11, 22, 10],\n[59, 13, 59, 12]]");
		$display("Expect: 59, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 4;
		pixel_array_in[0][2] = 61;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 43;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 17;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 13;
		pixel_array_in[2][3] = 56;
		pixel_array_in[3][0] = 57;
		pixel_array_in[3][1] = 3;
		pixel_array_in[3][2] = 22;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[5, 40, 52, 61],\n[44, 41, 54, 29],\n[14, 3, 45, 55],\n[7, 62, 29, 25]]");
		$display("Expect: 144, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 30;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 53;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 20;
		pixel_array_in[1][1] = 61;
		pixel_array_in[1][2] = 19;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 45;
		pixel_array_in[2][1] = 34;
		pixel_array_in[2][2] = 20;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 17;
		pixel_array_in[3][2] = 5;
		pixel_array_in[3][3] = 25;
		#10;
		
		$display("Input: \n[[19, 28, 34, 2],\n[25, 29, 62, 6],\n[30, 14, 51, 54],\n[25, 50, 36, 48]]");
		$display("Expect: 134, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 3;
		pixel_array_in[0][1] = 13;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 55;
		pixel_array_in[1][2] = 43;
		pixel_array_in[1][3] = 41;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 45;
		pixel_array_in[3][1] = 49;
		pixel_array_in[3][2] = 52;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[25, 5, 17, 55],\n[37, 44, 44, 48],\n[60, 38, 7, 23],\n[13, 15, 60, 54]]");
		$display("Expect: 177, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 60;
		pixel_array_in[1][0] = 30;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 59;
		pixel_array_in[2][0] = 41;
		pixel_array_in[2][1] = 46;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 6;
		pixel_array_in[3][0] = 20;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 51;
		#10;
		
		$display("Input: \n[[61, 4, 61, 12],\n[9, 27, 43, 48],\n[17, 38, 13, 56],\n[57, 3, 22, 44]]");
		$display("Expect: 135, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 26;
		pixel_array_in[0][1] = 3;
		pixel_array_in[0][2] = 40;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 10;
		pixel_array_in[1][2] = 26;
		pixel_array_in[1][3] = 14;
		pixel_array_in[2][0] = 18;
		pixel_array_in[2][1] = 31;
		pixel_array_in[2][2] = 33;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 30;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 5;
		#10;
		
		$display("Input: \n[[30, 19, 53, 44],\n[20, 61, 19, 25],\n[45, 34, 20, 39],\n[36, 17, 5, 25]]");
		$display("Expect: 210, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 35;
		pixel_array_in[0][1] = 53;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 38;
		pixel_array_in[1][0] = 55;
		pixel_array_in[1][1] = 44;
		pixel_array_in[1][2] = 45;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 20;
		pixel_array_in[2][1] = 8;
		pixel_array_in[2][2] = 11;
		pixel_array_in[2][3] = 20;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 9;
		#10;
		
		$display("Input: \n[[3, 13, 4, 57],\n[13, 55, 43, 41],\n[47, 12, 42, 53],\n[45, 49, 52, 33]]");
		$display("Expect: 198, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 43;
		pixel_array_in[0][1] = 34;
		pixel_array_in[0][2] = 29;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 49;
		pixel_array_in[1][1] = 51;
		pixel_array_in[1][2] = 49;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 29;
		pixel_array_in[3][2] = 19;
		pixel_array_in[3][3] = 45;
		#10;
		
		$display("Input: \n[[0, 40, 45, 60],\n[30, 35, 11, 59],\n[41, 46, 19, 6],\n[20, 50, 27, 51]]");
		$display("Expect: 122, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 7;
		pixel_array_in[0][1] = 15;
		pixel_array_in[0][2] = 15;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 55;
		pixel_array_in[1][2] = 23;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 24;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 62;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[26, 3, 40, 45],\n[13, 10, 26, 14],\n[18, 31, 33, 18],\n[30, 58, 3, 5]]");
		$display("Expect: 68, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 44;
		pixel_array_in[0][1] = 9;
		pixel_array_in[0][2] = 27;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 13;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 2;
		pixel_array_in[2][0] = 29;
		pixel_array_in[2][1] = 54;
		pixel_array_in[2][2] = 37;
		pixel_array_in[2][3] = 47;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 15;
		pixel_array_in[3][2] = 52;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[35, 53, 14, 38],\n[55, 44, 45, 0],\n[20, 8, 11, 20],\n[31, 32, 27, 9]]");
		$display("Expect: 145, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 59;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 27;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 58;
		pixel_array_in[2][1] = 6;
		pixel_array_in[2][2] = 37;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 10;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[43, 34, 29, 57],\n[49, 51, 49, 47],\n[31, 40, 30, 30],\n[29, 29, 19, 45]]");
		$display("Expect: 199, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 1;
		pixel_array_in[0][2] = 39;
		pixel_array_in[0][3] = 4;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 5;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 21;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 19;
		pixel_array_in[2][2] = 16;
		pixel_array_in[2][3] = 7;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 16;
		pixel_array_in[3][2] = 33;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[7, 15, 15, 0],\n[31, 55, 23, 56],\n[11, 24, 7, 30],\n[0, 18, 62, 7]]");
		$display("Expect: 183, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 14;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 43;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 19;
		pixel_array_in[2][0] = 36;
		pixel_array_in[2][1] = 6;
		pixel_array_in[2][2] = 28;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 2;
		pixel_array_in[3][2] = 18;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[44, 9, 27, 42],\n[9, 13, 22, 2],\n[29, 54, 37, 47],\n[61, 15, 52, 6]]");
		$display("Expect: 96, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 27;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 24;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 26;
		pixel_array_in[1][2] = 23;
		pixel_array_in[1][3] = 61;
		pixel_array_in[2][0] = 8;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 12;
		pixel_array_in[2][3] = 19;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 15;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 59;
		#10;
		
		$display("Input: \n[[19, 18, 59, 2],\n[27, 52, 39, 46],\n[58, 6, 37, 53],\n[23, 10, 12, 6]]");
		$display("Expect: 175, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 38;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 20;
		pixel_array_in[1][1] = 21;
		pixel_array_in[1][2] = 46;
		pixel_array_in[1][3] = 37;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 18;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 14;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 52;
		pixel_array_in[3][2] = 31;
		pixel_array_in[3][3] = 18;
		#10;
		
		$display("Input: \n[[8, 1, 39, 4],\n[38, 5, 37, 21],\n[50, 19, 16, 7],\n[46, 16, 33, 44]]");
		$display("Expect: 43, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 2;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 46;
		pixel_array_in[1][0] = 59;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 53;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 58;
		pixel_array_in[2][3] = 40;
		pixel_array_in[3][0] = 2;
		pixel_array_in[3][1] = 7;
		pixel_array_in[3][2] = 54;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[19, 14, 4, 59],\n[43, 25, 15, 19],\n[36, 6, 28, 3],\n[15, 2, 18, 60]]");
		$display("Expect: 79, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 48;
		pixel_array_in[0][1] = 16;
		pixel_array_in[0][2] = 5;
		pixel_array_in[0][3] = 5;
		pixel_array_in[1][0] = 55;
		pixel_array_in[1][1] = 38;
		pixel_array_in[1][2] = 44;
		pixel_array_in[1][3] = 58;
		pixel_array_in[2][0] = 49;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 56;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[27, 52, 24, 39],\n[61, 26, 23, 61],\n[8, 11, 12, 19],\n[31, 15, 7, 59]]");
		$display("Expect: 72, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 46;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 5;
		pixel_array_in[0][3] = 62;
		pixel_array_in[1][0] = 34;
		pixel_array_in[1][1] = 55;
		pixel_array_in[1][2] = 26;
		pixel_array_in[1][3] = 9;
		pixel_array_in[2][0] = 7;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 32;
		pixel_array_in[2][3] = 14;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 36;
		pixel_array_in[3][2] = 8;
		pixel_array_in[3][3] = 24;
		#10;
		
		$display("Input: \n[[53, 38, 51, 55],\n[20, 21, 46, 37],\n[47, 18, 57, 14],\n[40, 52, 31, 18]]");
		$display("Expect: 98, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 20;
		pixel_array_in[0][1] = 20;
		pixel_array_in[0][2] = 29;
		pixel_array_in[0][3] = 13;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 51;
		pixel_array_in[1][3] = 37;
		pixel_array_in[2][0] = 9;
		pixel_array_in[2][1] = 6;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 53;
		pixel_array_in[3][1] = 10;
		pixel_array_in[3][2] = 52;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[29, 2, 34, 46],\n[59, 45, 56, 56],\n[53, 11, 58, 40],\n[2, 7, 54, 2]]");
		$display("Expect: 173, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 55;
		pixel_array_in[0][1] = 57;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 52;
		pixel_array_in[1][0] = 60;
		pixel_array_in[1][1] = 17;
		pixel_array_in[1][2] = 24;
		pixel_array_in[1][3] = 8;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 27;
		pixel_array_in[2][3] = 28;
		pixel_array_in[3][0] = 62;
		pixel_array_in[3][1] = 5;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 13;
		#10;
		
		$display("Input: \n[[48, 16, 5, 5],\n[55, 38, 44, 58],\n[49, 35, 56, 10],\n[5, 57, 51, 44]]");
		$display("Expect: 158, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 20;
		pixel_array_in[0][1] = 21;
		pixel_array_in[0][2] = 25;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 55;
		pixel_array_in[1][1] = 21;
		pixel_array_in[1][2] = 16;
		pixel_array_in[1][3] = 61;
		pixel_array_in[2][0] = 46;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 26;
		pixel_array_in[3][0] = 14;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 23;
		#10;
		
		$display("Input: \n[[46, 52, 5, 62],\n[34, 55, 26, 9],\n[7, 38, 32, 14],\n[23, 36, 8, 24]]");
		$display("Expect: 197, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 31;
		pixel_array_in[0][1] = 3;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 22;
		pixel_array_in[1][0] = 19;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 51;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 55;
		pixel_array_in[2][3] = 50;
		pixel_array_in[3][0] = 56;
		pixel_array_in[3][1] = 47;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[20, 20, 29, 13],\n[44, 50, 51, 37],\n[9, 6, 5, 25],\n[53, 10, 52, 20]]");
		$display("Expect: 173, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 55;
		pixel_array_in[0][2] = 16;
		pixel_array_in[0][3] = 24;
		pixel_array_in[1][0] = 60;
		pixel_array_in[1][1] = 41;
		pixel_array_in[1][2] = 59;
		pixel_array_in[1][3] = 53;
		pixel_array_in[2][0] = 55;
		pixel_array_in[2][1] = 26;
		pixel_array_in[2][2] = 59;
		pixel_array_in[2][3] = 58;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 16;
		pixel_array_in[3][3] = 48;
		#10;
		
		$display("Input: \n[[55, 57, 21, 52],\n[60, 17, 24, 8],\n[11, 45, 27, 28],\n[62, 5, 48, 13]]");
		$display("Expect: 79, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 43;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 47;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 22;
		pixel_array_in[1][2] = 44;
		pixel_array_in[1][3] = 28;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 21;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 58;
		pixel_array_in[3][0] = 55;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 31;
		pixel_array_in[3][3] = 34;
		#10;
		
		$display("Input: \n[[20, 21, 25, 41],\n[55, 21, 16, 61],\n[46, 10, 62, 26],\n[14, 50, 15, 23]]");
		$display("Expect: 64, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 42;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 41;
		pixel_array_in[0][3] = 52;
		pixel_array_in[1][0] = 56;
		pixel_array_in[1][1] = 56;
		pixel_array_in[1][2] = 17;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 23;
		pixel_array_in[2][1] = 60;
		pixel_array_in[2][2] = 3;
		pixel_array_in[2][3] = 12;
		pixel_array_in[3][0] = 22;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 26;
		pixel_array_in[3][3] = 40;
		#10;
		
		$display("Input: \n[[31, 3, 21, 22],\n[19, 25, 51, 46],\n[0, 35, 55, 50],\n[56, 47, 32, 33]]");
		$display("Expect: 139, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 17;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 30;
		pixel_array_in[1][2] = 42;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 38;
		pixel_array_in[2][1] = 25;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 26;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 22;
		pixel_array_in[3][3] = 34;
		#10;
		
		$display("Input: \n[[53, 55, 16, 24],\n[60, 41, 59, 53],\n[55, 26, 59, 58],\n[40, 25, 16, 48]]");
		$display("Expect: 163, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 3;
		pixel_array_in[0][1] = 14;
		pixel_array_in[0][2] = 36;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 40;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 20;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 2;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 46;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[1, 43, 30, 47],\n[58, 22, 44, 28],\n[60, 21, 44, 58],\n[55, 18, 31, 34]]");
		$display("Expect: 90, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 44;
		pixel_array_in[0][1] = 9;
		pixel_array_in[0][2] = 37;
		pixel_array_in[0][3] = 16;
		pixel_array_in[1][0] = 52;
		pixel_array_in[1][1] = 6;
		pixel_array_in[1][2] = 38;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 18;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 19;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 41;
		#10;
		
		$display("Input: \n[[42, 25, 41, 52],\n[56, 56, 17, 17],\n[23, 60, 3, 12],\n[22, 45, 26, 40]]");
		$display("Expect: 201, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 47;
		pixel_array_in[0][1] = 13;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 2;
		pixel_array_in[1][1] = 39;
		pixel_array_in[1][2] = 31;
		pixel_array_in[1][3] = 50;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 48;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 8;
		#10;
		
		$display("Input: \n[[15, 58, 51, 17],\n[11, 30, 42, 4],\n[38, 25, 61, 26],\n[15, 30, 22, 34]]");
		$display("Expect: 129, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 43;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 14;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 59;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 1;
		pixel_array_in[3][3] = 10;
		#10;
		
		$display("Input: \n[[3, 14, 36, 10],\n[32, 40, 13, 47],\n[47, 20, 62, 24],\n[2, 13, 46, 12]]");
		$display("Expect: 136, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 34;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 17;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 30;
		pixel_array_in[2][2] = 21;
		pixel_array_in[2][3] = 2;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 53;
		#10;
		
		$display("Input: \n[[44, 9, 37, 16],\n[52, 6, 38, 29],\n[40, 18, 5, 19],\n[36, 28, 7, 41]]");
		$display("Expect: 39, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 46;
		pixel_array_in[0][3] = 7;
		pixel_array_in[1][0] = 23;
		pixel_array_in[1][1] = 39;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 38;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 60;
		pixel_array_in[2][3] = 17;
		pixel_array_in[3][0] = 60;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 13;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[47, 13, 32, 40],\n[2, 39, 31, 50],\n[12, 7, 62, 55],\n[48, 0, 59, 8]]");
		$display("Expect: 148, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 38;
		pixel_array_in[0][1] = 23;
		pixel_array_in[0][2] = 38;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 2;
		pixel_array_in[1][1] = 42;
		pixel_array_in[1][2] = 51;
		pixel_array_in[1][3] = 30;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 17;
		pixel_array_in[3][0] = 14;
		pixel_array_in[3][1] = 1;
		pixel_array_in[3][2] = 54;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[8, 45, 30, 1],\n[43, 23, 14, 39],\n[39, 59, 5, 36],\n[42, 30, 1, 10]]");
		$display("Expect: 96, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 33;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 35;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 52;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 8;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 37;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 1;
		pixel_array_in[3][2] = 30;
		pixel_array_in[3][3] = 17;
		#10;
		
		$display("Input: \n[[8, 34, 48, 10],\n[58, 0, 17, 48],\n[0, 30, 21, 2],\n[41, 59, 60, 53]]");
		$display("Expect: 6, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 56;
		pixel_array_in[0][1] = 12;
		pixel_array_in[0][2] = 3;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 44;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 52;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 34;
		pixel_array_in[2][2] = 8;
		pixel_array_in[2][3] = 20;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 62;
		pixel_array_in[3][2] = 19;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[21, 40, 46, 7],\n[23, 39, 30, 46],\n[38, 3, 60, 17],\n[60, 14, 13, 35]]");
		$display("Expect: 130, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 61;
		pixel_array_in[0][2] = 11;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 56;
		pixel_array_in[2][3] = 33;
		pixel_array_in[3][0] = 53;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 57;
		pixel_array_in[3][3] = 26;
		#10;
		
		$display("Input: \n[[38, 23, 38, 57],\n[2, 42, 51, 30],\n[47, 57, 30, 17],\n[14, 1, 54, 52]]");
		$display("Expect: 203, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 62;
		pixel_array_in[0][2] = 40;
		pixel_array_in[0][3] = 20;
		pixel_array_in[1][0] = 51;
		pixel_array_in[1][1] = 53;
		pixel_array_in[1][2] = 58;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 56;
		pixel_array_in[2][1] = 41;
		pixel_array_in[2][2] = 26;
		pixel_array_in[2][3] = 23;
		pixel_array_in[3][0] = 14;
		pixel_array_in[3][1] = 53;
		pixel_array_in[3][2] = 28;
		pixel_array_in[3][3] = 31;
		#10;
		
		$display("Input: \n[[33, 56, 14, 36],\n[35, 37, 52, 12],\n[8, 10, 37, 36],\n[42, 1, 30, 17]]");
		$display("Expect: 142, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 4;
		pixel_array_in[0][1] = 27;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 39;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 50;
		pixel_array_in[2][0] = 33;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 26;
		pixel_array_in[2][3] = 19;
		pixel_array_in[3][0] = 51;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[56, 12, 3, 1],\n[0, 44, 25, 52],\n[30, 34, 8, 20],\n[5, 62, 19, 33]]");
		$display("Expect: 167, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 55;
		pixel_array_in[0][1] = 27;
		pixel_array_in[0][2] = 10;
		pixel_array_in[0][3] = 37;
		pixel_array_in[1][0] = 7;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 47;
		pixel_array_in[1][3] = 30;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 18;
		pixel_array_in[2][2] = 16;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 53;
		#10;
		
		$display("Input: \n[[8, 61, 11, 19],\n[28, 28, 33, 6],\n[22, 45, 56, 33],\n[53, 44, 57, 26]]");
		$display("Expect: 127, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 11;
		pixel_array_in[0][1] = 24;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 15;
		pixel_array_in[1][2] = 16;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 14;
		pixel_array_in[3][0] = 16;
		pixel_array_in[3][1] = 53;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[1, 62, 40, 20],\n[51, 53, 58, 38],\n[56, 41, 26, 23],\n[14, 53, 28, 31]]");
		$display("Expect: 201, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 27;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 60;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 34;
		pixel_array_in[2][1] = 14;
		pixel_array_in[2][2] = 6;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 27;
		pixel_array_in[3][1] = 40;
		pixel_array_in[3][2] = 8;
		pixel_array_in[3][3] = 22;
		#10;
		
		$display("Input: \n[[4, 27, 30, 36],\n[61, 39, 11, 50],\n[33, 11, 26, 19],\n[51, 42, 29, 35]]");
		$display("Expect: 106, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 14;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 48;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 20;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 24;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 19;
		pixel_array_in[3][0] = 2;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 62;
		pixel_array_in[3][3] = 47;
		#10;
		
		$display("Input: \n[[55, 27, 10, 37],\n[7, 1, 47, 30],\n[42, 18, 16, 49],\n[41, 18, 6, 53]]");
		$display("Expect: 42, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 60;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 30;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 9;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 56;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 51;
		pixel_array_in[3][0] = 21;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[11, 24, 51, 10],\n[11, 15, 16, 25],\n[1, 45, 17, 14],\n[16, 53, 59, 1]]");
		$display("Expect: 77, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 55;
		pixel_array_in[0][1] = 33;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 35;
		pixel_array_in[1][0] = 41;
		pixel_array_in[1][1] = 39;
		pixel_array_in[1][2] = 55;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 53;
		pixel_array_in[2][3] = 23;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 3;
		#10;
		
		$display("Input: \n[[27, 54, 45, 1],\n[60, 32, 10, 62],\n[34, 14, 6, 24],\n[27, 40, 8, 22]]");
		$display("Expect: 75, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 11;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 57;
		pixel_array_in[0][3] = 61;
		pixel_array_in[1][0] = 41;
		pixel_array_in[1][1] = 44;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 33;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 31;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 28;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[61, 14, 51, 48],\n[10, 49, 20, 6],\n[12, 24, 23, 19],\n[2, 44, 62, 47]]");
		$display("Expect: 172, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 13;
		pixel_array_in[0][1] = 62;
		pixel_array_in[0][2] = 36;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 9;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 28;
		pixel_array_in[2][0] = 9;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 3;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 49;
		pixel_array_in[3][1] = 53;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Input: \n[[57, 60, 23, 45],\n[11, 30, 25, 9],\n[10, 56, 57, 51],\n[21, 13, 29, 56]]");
		$display("Expect: 144, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 53;
		pixel_array_in[0][2] = 1;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 16;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[55, 33, 21, 35],\n[41, 39, 55, 29],\n[31, 55, 53, 23],\n[23, 13, 59, 3]]");
		$display("Expect: 189, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[11, 10, 57, 61],\n[41, 44, 36, 33],\n[60, 3, 31, 3],\n[32, 48, 28, 35]]");
		$display("Expect: 142, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[13, 62, 36, 33],\n[0, 9, 50, 28],\n[9, 40, 3, 44],\n[49, 53, 6, 0]]");
		$display("Expect: 73, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[21, 53, 1, 53],\n[32, 12, 5, 32],\n[24, 10, 57, 32],\n[40, 59, 16, 56]]");
		$display("Expect: 29, Result: %d", pixel_out);
		$display("");
		#10;
		
		
		$display("Finishing Sim"); //print nice message
		$finish;
		
    end
endmodule //counter_tb

`default_nettype wire