`timescale 1ns / 1ps
`default_nettype none

module kernel_1_tb;

    //make logics for inputs and outputs!
    logic clk_in;
    logic rst_in;
    logic valid_in;
    logic [5:0] pixel_array_in [3:0][3:0];
    logic [8:0] pixel_out;

    kernel_1 uut (
        .clk_in(clk_in),
        .p1(pixel_array_in[0][1]),
        .p2(pixel_array_in[1][1]),
        .p3(pixel_array_in[2][1]),
        .p4(pixel_array_in[3][1]),
        .pixel_out(pixel_out)
    );
    always begin
        #5;  //every 5 ns switch...so period of clock is 10 ns...100 MHz clock
        clk_in = !clk_in;
    end

    //initial block...this is our test simulation
    initial begin
        
		$dumpfile("test/kernel_1.vcd"); //file to store value change dump (vcd)
		$dumpvars(0,kernel_1_tb); //store everything at the current level and below
		$display("Starting Sim"); //print nice message
		clk_in = 0; //initialize clk (super important)
		rst_in = 0; //initialize rst (super important)
		
		#10;  //wait a little bit of time at beginning
		rst_in = 1; //reset system
		#10; //hold high for a few clock cycles
		rst_in=0;
		
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 0;
		#10;
		
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 32;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 32;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 32;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 32;
		#10;
		
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 63;
		#10;
		
		$display("Input: \n[[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0]]");
		$display("Expect: 0, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 63;
		#10;
		
		$display("Input: \n[[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32]]");
		$display("Expect: 128, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Input: \n[[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63]]");
		$display("Expect: 252, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 38;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 1;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 35;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 34;
		pixel_array_in[2][3] = 61;
		pixel_array_in[3][0] = 37;
		pixel_array_in[3][1] = 47;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 57;
		#10;
		
		$display("Input: \n[[63, 0, 0, 63],\n[0, 63, 63, 0],\n[0, 63, 63, 0],\n[63, 0, 0, 63]]");
		$display("Expect: 384>val>255, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 47;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 57;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 26;
		pixel_array_in[1][2] = 58;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 59;
		pixel_array_in[2][1] = 61;
		pixel_array_in[2][2] = 21;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 43;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 42;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[0, 63, 63, 0],\n[63, 0, 0, 63],\n[63, 0, 0, 63],\n[0, 63, 63, 0]]");
		$display("Expect: val>383, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 51;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 18;
		pixel_array_in[1][2] = 14;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 35;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 60;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 25;
		#10;
		
		$display("Input: \n[[15, 18, 38, 1],\n[1, 32, 30, 39],\n[35, 3, 34, 61],\n[37, 47, 42, 57]]");
		$display("Expect: 104, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 6;
		pixel_array_in[1][0] = 23;
		pixel_array_in[1][1] = 59;
		pixel_array_in[1][2] = 4;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 46;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 17;
		pixel_array_in[3][2] = 5;
		pixel_array_in[3][3] = 41;
		#10;
		
		$display("Input: \n[[47, 48, 57, 55],\n[58, 26, 58, 62],\n[59, 61, 21, 32],\n[43, 59, 42, 27]]");
		$display("Expect: 126, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 34;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 14;
		pixel_array_in[1][2] = 18;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 19;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 9;
		pixel_array_in[2][3] = 7;
		pixel_array_in[3][0] = 60;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 41;
		pixel_array_in[3][3] = 19;
		#10;
		
		$display("Input: \n[[51, 25, 52, 10],\n[9, 18, 14, 0],\n[42, 35, 35, 1],\n[60, 57, 2, 25]]");
		$display("Expect: 81, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 47;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 28;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 47;
		pixel_array_in[1][2] = 34;
		pixel_array_in[1][3] = 61;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 38;
		pixel_array_in[3][0] = 39;
		pixel_array_in[3][1] = 4;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 5;
		#10;
		
		$display("Input: \n[[25, 40, 51, 6],\n[23, 59, 4, 12],\n[0, 3, 61, 46],\n[13, 17, 5, 41]]");
		$display("Expect: 194, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 45;
		pixel_array_in[0][1] = 38;
		pixel_array_in[0][2] = 36;
		pixel_array_in[0][3] = 37;
		pixel_array_in[1][0] = 20;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 53;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 55;
		pixel_array_in[2][1] = 24;
		pixel_array_in[2][2] = 2;
		pixel_array_in[2][3] = 5;
		pixel_array_in[3][0] = 33;
		pixel_array_in[3][1] = 53;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[61, 45, 34, 34],\n[61, 14, 18, 32],\n[19, 40, 9, 7],\n[60, 0, 41, 19]]");
		$display("Expect: 72, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 22;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 3;
		pixel_array_in[1][1] = 62;
		pixel_array_in[1][2] = 2;
		pixel_array_in[1][3] = 53;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 50;
		pixel_array_in[2][2] = 18;
		pixel_array_in[2][3] = 35;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[47, 56, 7, 28],\n[10, 47, 34, 61],\n[24, 11, 52, 38],\n[39, 4, 55, 5]]");
		$display("Expect: 156, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 44;
		pixel_array_in[0][1] = 36;
		pixel_array_in[0][2] = 33;
		pixel_array_in[0][3] = 20;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 55;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 2;
		pixel_array_in[2][0] = 41;
		pixel_array_in[2][1] = 25;
		pixel_array_in[2][2] = 12;
		pixel_array_in[2][3] = 26;
		pixel_array_in[3][0] = 48;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[45, 38, 36, 37],\n[20, 1, 53, 35],\n[55, 24, 2, 5],\n[33, 53, 17, 56]]");
		$display("Expect: 9, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 33;
		pixel_array_in[0][1] = 27;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 27;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 12;
		pixel_array_in[1][3] = 53;
		pixel_array_in[2][0] = 18;
		pixel_array_in[2][1] = 58;
		pixel_array_in[2][2] = 31;
		pixel_array_in[2][3] = 46;
		pixel_array_in[3][0] = 20;
		pixel_array_in[3][1] = 8;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 23;
		#10;
		
		$display("Input: \n[[21, 10, 22, 12],\n[3, 62, 2, 53],\n[42, 50, 18, 35],\n[0, 30, 12, 27]]");
		$display("Expect: 254, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 49;
		pixel_array_in[0][1] = 24;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 30;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 55;
		pixel_array_in[1][3] = 41;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 20;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 37;
		pixel_array_in[3][1] = 35;
		pixel_array_in[3][2] = 25;
		pixel_array_in[3][3] = 15;
		#10;
		
		$display("Input: \n[[44, 36, 33, 20],\n[58, 55, 33, 2],\n[41, 25, 12, 26],\n[48, 57, 3, 1]]");
		$display("Expect: 197, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 53;
		pixel_array_in[0][2] = 40;
		pixel_array_in[0][3] = 16;
		pixel_array_in[1][0] = 20;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 15;
		pixel_array_in[2][2] = 35;
		pixel_array_in[2][3] = 4;
		pixel_array_in[3][0] = 39;
		pixel_array_in[3][1] = 24;
		pixel_array_in[3][2] = 35;
		pixel_array_in[3][3] = 23;
		#10;
		
		$display("Input: \n[[33, 27, 12, 44],\n[27, 7, 12, 53],\n[18, 58, 31, 46],\n[20, 8, 7, 23]]");
		$display("Expect: 68, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 49;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 20;
		pixel_array_in[1][1] = 42;
		pixel_array_in[1][2] = 46;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 46;
		pixel_array_in[2][2] = 2;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 55;
		pixel_array_in[3][1] = 29;
		pixel_array_in[3][2] = 10;
		pixel_array_in[3][3] = 32;
		#10;
		
		$display("Input: \n[[49, 24, 32, 30],\n[22, 50, 55, 41],\n[24, 20, 54, 55],\n[37, 35, 25, 15]]");
		$display("Expect: 181, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 14;
		pixel_array_in[0][1] = 37;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 9;
		pixel_array_in[2][1] = 42;
		pixel_array_in[2][2] = 14;
		pixel_array_in[2][3] = 52;
		pixel_array_in[3][0] = 24;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 33;
		pixel_array_in[3][3] = 21;
		#10;
		
		$display("Input: \n[[32, 53, 40, 16],\n[20, 35, 15, 17],\n[40, 15, 35, 4],\n[39, 24, 35, 23]]");
		$display("Expect: 117, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 62;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 61;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 47;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 51;
		pixel_array_in[2][2] = 38;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 57;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 43;
		#10;
		
		$display("Input: \n[[49, 54, 7, 10],\n[20, 42, 46, 39],\n[0, 46, 2, 9],\n[55, 29, 10, 32]]");
		$display("Expect: 169, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 45;
		pixel_array_in[0][1] = 8;
		pixel_array_in[0][2] = 49;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 58;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 62;
		pixel_array_in[2][1] = 60;
		pixel_array_in[2][2] = 21;
		pixel_array_in[2][3] = 4;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 16;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 43;
		#10;
		
		$display("Input: \n[[14, 37, 21, 18],\n[13, 45, 50, 62],\n[9, 42, 14, 52],\n[24, 26, 33, 21]]");
		$display("Expect: 181, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 50;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 5;
		pixel_array_in[0][3] = 50;
		pixel_array_in[1][0] = 35;
		pixel_array_in[1][1] = 39;
		pixel_array_in[1][2] = 12;
		pixel_array_in[1][3] = 60;
		pixel_array_in[2][0] = 56;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 13;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 20;
		pixel_array_in[3][1] = 47;
		pixel_array_in[3][2] = 16;
		pixel_array_in[3][3] = 14;
		#10;
		
		$display("Input: \n[[0, 62, 48, 61],\n[57, 12, 47, 4],\n[12, 51, 38, 36],\n[57, 13, 12, 43]]");
		$display("Expect: 69, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 36;
		pixel_array_in[0][1] = 60;
		pixel_array_in[0][2] = 57;
		pixel_array_in[0][3] = 4;
		pixel_array_in[1][0] = 2;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 58;
		pixel_array_in[3][0] = 43;
		pixel_array_in[3][1] = 40;
		pixel_array_in[3][2] = 9;
		pixel_array_in[3][3] = 61;
		#10;
		
		$display("Input: \n[[45, 8, 49, 2],\n[57, 58, 33, 17],\n[62, 60, 21, 4],\n[0, 16, 59, 43]]");
		$display("Expect: 251, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 34;
		pixel_array_in[0][1] = 6;
		pixel_array_in[0][2] = 50;
		pixel_array_in[0][3] = 47;
		pixel_array_in[1][0] = 50;
		pixel_array_in[1][1] = 15;
		pixel_array_in[1][2] = 48;
		pixel_array_in[1][3] = 22;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 48;
		pixel_array_in[2][2] = 12;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 8;
		pixel_array_in[3][1] = 24;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 41;
		#10;
		
		$display("Input: \n[[50, 54, 5, 50],\n[35, 39, 12, 60],\n[56, 55, 13, 0],\n[20, 47, 16, 14]]");
		$display("Expect: 165, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 14;
		pixel_array_in[0][1] = 6;
		pixel_array_in[0][2] = 43;
		pixel_array_in[0][3] = 44;
		pixel_array_in[1][0] = 10;
		pixel_array_in[1][1] = 13;
		pixel_array_in[1][2] = 62;
		pixel_array_in[1][3] = 33;
		pixel_array_in[2][0] = 46;
		pixel_array_in[2][1] = 2;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 53;
		pixel_array_in[3][1] = 4;
		pixel_array_in[3][2] = 28;
		pixel_array_in[3][3] = 37;
		#10;
		
		$display("Input: \n[[36, 60, 57, 4],\n[2, 49, 30, 35],\n[50, 12, 23, 58],\n[43, 40, 9, 61]]");
		$display("Expect: 160, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 20;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 43;
		pixel_array_in[0][3] = 46;
		pixel_array_in[1][0] = 21;
		pixel_array_in[1][1] = 62;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 14;
		pixel_array_in[2][0] = 52;
		pixel_array_in[2][1] = 6;
		pixel_array_in[2][2] = 27;
		pixel_array_in[2][3] = 46;
		pixel_array_in[3][0] = 56;
		pixel_array_in[3][1] = 2;
		pixel_array_in[3][2] = 35;
		pixel_array_in[3][3] = 45;
		#10;
		
		$display("Input: \n[[34, 6, 50, 47],\n[50, 15, 48, 22],\n[40, 48, 12, 43],\n[8, 24, 55, 41]]");
		$display("Expect: 91, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 50;
		pixel_array_in[0][1] = 11;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 3;
		pixel_array_in[1][1] = 39;
		pixel_array_in[1][2] = 42;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 28;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 1;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 40;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[14, 6, 43, 44],\n[10, 13, 62, 33],\n[46, 2, 19, 44],\n[53, 4, 28, 37]]");
		$display("Expect: 44, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 59;
		pixel_array_in[0][2] = 62;
		pixel_array_in[0][3] = 23;
		pixel_array_in[1][0] = 19;
		pixel_array_in[1][1] = 51;
		pixel_array_in[1][2] = 38;
		pixel_array_in[1][3] = 26;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 23;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 25;
		pixel_array_in[3][3] = 30;
		#10;
		
		$display("Input: \n[[20, 40, 43, 46],\n[21, 62, 11, 14],\n[52, 6, 27, 46],\n[56, 2, 35, 45]]");
		$display("Expect: 209, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 54;
		pixel_array_in[0][3] = 56;
		pixel_array_in[1][0] = 30;
		pixel_array_in[1][1] = 30;
		pixel_array_in[1][2] = 59;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 45;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 21;
		pixel_array_in[3][0] = 6;
		pixel_array_in[3][1] = 19;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 34;
		#10;
		
		$display("Input: \n[[50, 11, 21, 59],\n[3, 39, 42, 12],\n[28, 36, 52, 62],\n[1, 57, 40, 33]]");
		$display("Expect: 159, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 11;
		pixel_array_in[0][1] = 35;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 23;
		pixel_array_in[1][0] = 40;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 31;
		pixel_array_in[1][3] = 40;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 22;
		pixel_array_in[3][1] = 9;
		pixel_array_in[3][2] = 52;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[32, 59, 62, 23],\n[19, 51, 38, 26],\n[15, 23, 19, 23],\n[10, 58, 25, 30]]");
		$display("Expect: 175, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 59;
		pixel_array_in[0][1] = 44;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 47;
		pixel_array_in[1][0] = 30;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 44;
		pixel_array_in[1][3] = 16;
		pixel_array_in[2][0] = 2;
		pixel_array_in[2][1] = 28;
		pixel_array_in[2][2] = 13;
		pixel_array_in[2][3] = 27;
		pixel_array_in[3][0] = 16;
		pixel_array_in[3][1] = 22;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 48;
		#10;
		
		$display("Input: \n[[22, 40, 54, 56],\n[30, 30, 59, 46],\n[45, 10, 43, 21],\n[6, 19, 17, 34]]");
		$display("Expect: 100, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 56;
		pixel_array_in[0][1] = 4;
		pixel_array_in[0][2] = 59;
		pixel_array_in[0][3] = 16;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 57;
		pixel_array_in[1][3] = 62;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 60;
		pixel_array_in[3][1] = 52;
		pixel_array_in[3][2] = 49;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[11, 35, 52, 23],\n[40, 33, 31, 40],\n[40, 44, 57, 3],\n[22, 9, 52, 2]]");
		$display("Expect: 143, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 23;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 17;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 62;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 21;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 43;
		pixel_array_in[3][2] = 39;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[59, 44, 55, 47],\n[30, 23, 44, 16],\n[2, 28, 13, 27],\n[16, 22, 61, 48]]");
		$display("Expect: 90, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 23;
		pixel_array_in[0][1] = 47;
		pixel_array_in[0][2] = 6;
		pixel_array_in[0][3] = 51;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 38;
		pixel_array_in[1][2] = 7;
		pixel_array_in[1][3] = 1;
		pixel_array_in[2][0] = 3;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 24;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 31;
		pixel_array_in[3][2] = 53;
		pixel_array_in[3][3] = 57;
		#10;
		
		$display("Input: \n[[56, 4, 59, 16],\n[47, 52, 57, 62],\n[47, 11, 5, 30],\n[60, 52, 49, 16]]");
		$display("Expect: 184, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 22;
		pixel_array_in[0][2] = 5;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 50;
		pixel_array_in[1][1] = 41;
		pixel_array_in[1][2] = 24;
		pixel_array_in[1][3] = 49;
		pixel_array_in[2][0] = 16;
		pixel_array_in[2][1] = 52;
		pixel_array_in[2][2] = 6;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 40;
		pixel_array_in[3][1] = 19;
		pixel_array_in[3][2] = 19;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[23, 48, 17, 33],\n[62, 45, 13, 0],\n[21, 23, 19, 62],\n[5, 43, 39, 12]]");
		$display("Expect: 159, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 31;
		pixel_array_in[0][2] = 60;
		pixel_array_in[0][3] = 23;
		pixel_array_in[1][0] = 24;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 53;
		pixel_array_in[1][3] = 11;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 54;
		pixel_array_in[2][2] = 27;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 44;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 21;
		#10;
		
		$display("Input: \n[[23, 47, 6, 51],\n[57, 38, 7, 1],\n[3, 57, 24, 43],\n[17, 31, 53, 57]]");
		$display("Expect: 167, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 52;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 8;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 52;
		pixel_array_in[1][1] = 38;
		pixel_array_in[1][2] = 60;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 37;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 27;
		pixel_array_in[3][2] = 47;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[57, 22, 5, 19],\n[50, 41, 24, 49],\n[16, 52, 6, 43],\n[40, 19, 19, 20]]");
		$display("Expect: 181, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 1;
		pixel_array_in[0][2] = 39;
		pixel_array_in[0][3] = 23;
		pixel_array_in[1][0] = 39;
		pixel_array_in[1][1] = 4;
		pixel_array_in[1][2] = 60;
		pixel_array_in[1][3] = 55;
		pixel_array_in[2][0] = 61;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 4;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 39;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[15, 31, 60, 23],\n[24, 52, 53, 11],\n[57, 54, 27, 53],\n[44, 30, 56, 21]]");
		$display("Expect: 217, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 6;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 1;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 42;
		pixel_array_in[1][1] = 1;
		pixel_array_in[1][2] = 48;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 58;
		pixel_array_in[2][1] = 4;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 47;
		pixel_array_in[3][3] = 46;
		#10;
		
		$display("Input: \n[[52, 56, 8, 12],\n[52, 38, 60, 15],\n[10, 37, 52, 32],\n[42, 27, 47, 27]]");
		$display("Expect: 147, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 37;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 61;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 9;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 43;
		pixel_array_in[2][0] = 25;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 51;
		pixel_array_in[2][3] = 16;
		pixel_array_in[3][0] = 34;
		pixel_array_in[3][1] = 41;
		pixel_array_in[3][2] = 18;
		pixel_array_in[3][3] = 5;
		#10;
		
		$display("Input: \n[[8, 1, 39, 23],\n[39, 4, 60, 55],\n[61, 35, 4, 0],\n[5, 45, 39, 58]]");
		$display("Expect: 41, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 58;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 26;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 36;
		pixel_array_in[1][1] = 31;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 16;
		pixel_array_in[2][0] = 53;
		pixel_array_in[2][1] = 6;
		pixel_array_in[2][2] = 37;
		pixel_array_in[2][3] = 33;
		pixel_array_in[3][0] = 28;
		pixel_array_in[3][1] = 11;
		pixel_array_in[3][2] = 38;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[6, 40, 1, 10],\n[42, 1, 48, 38],\n[58, 4, 22, 10],\n[46, 18, 47, 46]]");
		$display("Expect: val>383, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 5;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 30;
		pixel_array_in[1][0] = 25;
		pixel_array_in[1][1] = 56;
		pixel_array_in[1][2] = 40;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 36;
		pixel_array_in[2][3] = 22;
		pixel_array_in[3][0] = 44;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 62;
		#10;
		
		$display("Input: \n[[37, 56, 0, 61],\n[57, 9, 36, 43],\n[25, 55, 51, 16],\n[34, 41, 18, 5]]");
		$display("Expect: 61, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 34;
		pixel_array_in[0][1] = 1;
		pixel_array_in[0][2] = 18;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 15;
		pixel_array_in[1][1] = 59;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 54;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 25;
		pixel_array_in[2][2] = 11;
		pixel_array_in[2][3] = 11;
		pixel_array_in[3][0] = 34;
		pixel_array_in[3][1] = 10;
		pixel_array_in[3][2] = 57;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[58, 28, 26, 40],\n[36, 31, 33, 16],\n[53, 6, 37, 33],\n[28, 11, 38, 39]]");
		$display("Expect: 104, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 30;
		pixel_array_in[0][1] = 37;
		pixel_array_in[0][2] = 62;
		pixel_array_in[0][3] = 49;
		pixel_array_in[1][0] = 51;
		pixel_array_in[1][1] = 51;
		pixel_array_in[1][2] = 44;
		pixel_array_in[1][3] = 6;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 37;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 21;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 25;
		#10;
		
		$display("Input: \n[[15, 5, 45, 30],\n[25, 56, 40, 46],\n[31, 55, 36, 22],\n[44, 32, 45, 62]]");
		$display("Expect: 239, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 24;
		pixel_array_in[0][1] = 51;
		pixel_array_in[0][2] = 41;
		pixel_array_in[0][3] = 29;
		pixel_array_in[1][0] = 50;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 55;
		pixel_array_in[2][3] = 46;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 39;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[34, 1, 18, 40],\n[15, 59, 25, 54],\n[10, 25, 11, 11],\n[34, 10, 57, 52]]");
		$display("Expect: 226, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 3;
		pixel_array_in[0][1] = 29;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 13;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 9;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 58;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 13;
		pixel_array_in[3][0] = 57;
		pixel_array_in[3][1] = 7;
		pixel_array_in[3][2] = 54;
		pixel_array_in[3][3] = 43;
		#10;
		
		$display("Input: \n[[30, 37, 62, 49],\n[51, 51, 44, 6],\n[1, 37, 49, 36],\n[21, 55, 61, 25]]");
		$display("Expect: 194, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 2;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 30;
		pixel_array_in[1][3] = 26;
		pixel_array_in[2][0] = 33;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 44;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 55;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[24, 51, 41, 29],\n[50, 28, 0, 25],\n[47, 1, 55, 46],\n[5, 39, 59, 2]]");
		$display("Expect: 80, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 41;
		pixel_array_in[0][2] = 2;
		pixel_array_in[0][3] = 38;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 40;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 49;
		pixel_array_in[2][0] = 18;
		pixel_array_in[2][1] = 34;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 60;
		pixel_array_in[3][2] = 46;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[3, 29, 14, 2],\n[0, 13, 36, 9],\n[15, 58, 47, 13],\n[57, 7, 54, 43]]");
		$display("Expect: 88, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 54;
		pixel_array_in[0][1] = 16;
		pixel_array_in[0][2] = 51;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 48;
		pixel_array_in[1][1] = 57;
		pixel_array_in[1][2] = 14;
		pixel_array_in[1][3] = 57;
		pixel_array_in[2][0] = 41;
		pixel_array_in[2][1] = 43;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 37;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 43;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 31;
		#10;
		
		$display("Input: \n[[9, 2, 52, 40],\n[46, 35, 30, 26],\n[33, 36, 23, 53],\n[44, 37, 55, 44]]");
		$display("Expect: 150, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 41;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 8;
		pixel_array_in[0][3] = 3;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 22;
		pixel_array_in[1][2] = 52;
		pixel_array_in[1][3] = 30;
		pixel_array_in[2][0] = 53;
		pixel_array_in[2][1] = 56;
		pixel_array_in[2][2] = 14;
		pixel_array_in[2][3] = 38;
		pixel_array_in[3][0] = 54;
		pixel_array_in[3][1] = 7;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[22, 41, 2, 38],\n[11, 40, 3, 49],\n[18, 34, 22, 25],\n[31, 60, 46, 52]]");
		$display("Expect: 152, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 41;
		pixel_array_in[0][1] = 21;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 5;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 21;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 27;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 11;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 44;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 14;
		pixel_array_in[3][3] = 36;
		#10;
		
		$display("Input: \n[[54, 16, 51, 57],\n[48, 57, 14, 57],\n[41, 43, 62, 37],\n[31, 43, 15, 31]]");
		$display("Expect: 228, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 27;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 27;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 2;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 25;
		pixel_array_in[2][3] = 45;
		pixel_array_in[3][0] = 53;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 8;
		#10;
		
		$display("Input: \n[[41, 28, 8, 3],\n[13, 22, 52, 30],\n[53, 56, 14, 38],\n[54, 7, 7, 42]]");
		$display("Expect: 118, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 62;
		pixel_array_in[0][1] = 34;
		pixel_array_in[0][2] = 54;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 39;
		pixel_array_in[1][1] = 17;
		pixel_array_in[1][2] = 54;
		pixel_array_in[1][3] = 24;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 31;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 24;
		pixel_array_in[3][3] = 14;
		#10;
		
		$display("Input: \n[[41, 21, 30, 5],\n[61, 21, 32, 17],\n[27, 1, 11, 36],\n[44, 59, 14, 36]]");
		$display("Expect: 62, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 55;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 20;
		pixel_array_in[1][1] = 14;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 25;
		pixel_array_in[2][0] = 18;
		pixel_array_in[2][1] = 5;
		pixel_array_in[2][2] = 35;
		pixel_array_in[2][3] = 38;
		pixel_array_in[3][0] = 59;
		pixel_array_in[3][1] = 52;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 62;
		#10;
		
		$display("Input: \n[[22, 27, 55, 27],\n[57, 25, 37, 2],\n[11, 23, 25, 45],\n[53, 26, 12, 8]]");
		$display("Expect: 97, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 62;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 1;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 36;
		pixel_array_in[1][1] = 22;
		pixel_array_in[1][2] = 20;
		pixel_array_in[1][3] = 40;
		pixel_array_in[2][0] = 13;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 58;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[62, 34, 54, 18],\n[39, 17, 54, 24],\n[30, 32, 31, 62],\n[36, 32, 24, 14]]");
		$display("Expect: 75, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 2;
		pixel_array_in[0][3] = 3;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 4;
		pixel_array_in[1][2] = 28;
		pixel_array_in[1][3] = 16;
		pixel_array_in[2][0] = 2;
		pixel_array_in[2][1] = 53;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 11;
		pixel_array_in[3][1] = 54;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[53, 55, 23, 58],\n[20, 14, 33, 25],\n[18, 5, 35, 38],\n[59, 52, 17, 62]]");
		$display("Expect: 32, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 46;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 49;
		pixel_array_in[1][0] = 1;
		pixel_array_in[1][1] = 29;
		pixel_array_in[1][2] = 55;
		pixel_array_in[1][3] = 43;
		pixel_array_in[2][0] = 56;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 2;
		pixel_array_in[2][3] = 21;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 1;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 22;
		#10;
		
		$display("Input: \n[[62, 54, 1, 19],\n[36, 22, 20, 40],\n[13, 32, 47, 49],\n[38, 42, 58, 12]]");
		$display("Expect: 86, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 9;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 61;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 62;
		pixel_array_in[2][1] = 42;
		pixel_array_in[2][2] = 59;
		pixel_array_in[2][3] = 35;
		pixel_array_in[3][0] = 43;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 49;
		#10;
		
		$display("Input: \n[[1, 25, 2, 3],\n[47, 4, 28, 16],\n[2, 53, 52, 24],\n[11, 54, 48, 6]]");
		$display("Expect: 49, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 42;
		pixel_array_in[0][1] = 57;
		pixel_array_in[0][2] = 43;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 40;
		pixel_array_in[1][1] = 57;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 60;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 45;
		pixel_array_in[2][2] = 4;
		pixel_array_in[2][3] = 4;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 2;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 49;
		#10;
		
		$display("Input: \n[[46, 40, 45, 49],\n[1, 29, 55, 43],\n[56, 38, 2, 21],\n[19, 1, 32, 22]]");
		$display("Expect: 123, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 42;
		pixel_array_in[0][1] = 49;
		pixel_array_in[0][2] = 1;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 37;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 43;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 50;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 23;
		pixel_array_in[3][2] = 16;
		pixel_array_in[3][3] = 19;
		#10;
		
		$display("Input: \n[[29, 48, 55, 9],\n[11, 33, 61, 44],\n[62, 42, 59, 35],\n[43, 26, 61, 49]]");
		$display("Expect: 136, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 57;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 7;
		pixel_array_in[1][1] = 17;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 14;
		pixel_array_in[2][0] = 20;
		pixel_array_in[2][1] = 48;
		pixel_array_in[2][2] = 20;
		pixel_array_in[2][3] = 13;
		pixel_array_in[3][0] = 22;
		pixel_array_in[3][1] = 15;
		pixel_array_in[3][2] = 26;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[42, 57, 43, 19],\n[40, 57, 10, 60],\n[42, 45, 4, 4],\n[46, 2, 6, 49]]");
		$display("Expect: 222, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 55;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 62;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 45;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 24;
		pixel_array_in[1][3] = 5;
		pixel_array_in[2][0] = 3;
		pixel_array_in[2][1] = 42;
		pixel_array_in[2][2] = 58;
		pixel_array_in[2][3] = 57;
		pixel_array_in[3][0] = 26;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Input: \n[[42, 49, 1, 40],\n[37, 35, 43, 35],\n[39, 1, 50, 9],\n[15, 23, 16, 19]]");
		$display("Expect: 106, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 40;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 56;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 6;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 2;
		pixel_array_in[2][1] = 56;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 31;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 45;
		#10;
		
		$display("Input: \n[[57, 57, 34, 58],\n[7, 17, 10, 14],\n[20, 48, 20, 13],\n[22, 15, 26, 12]]");
		$display("Expect: 85, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 27;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 61;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 6;
		pixel_array_in[1][2] = 49;
		pixel_array_in[1][3] = 45;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 27;
		pixel_array_in[2][2] = 2;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 60;
		pixel_array_in[3][2] = 22;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[55, 17, 62, 10],\n[45, 28, 24, 5],\n[3, 42, 58, 57],\n[26, 44, 56, 0]]");
		$display("Expect: 126, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 30;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 39;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 29;
		pixel_array_in[1][1] = 11;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 57;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 53;
		pixel_array_in[2][2] = 58;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 27;
		pixel_array_in[3][1] = 22;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 23;
		#10;
		
		$display("Input: \n[[1, 40, 55, 56],\n[44, 35, 6, 48],\n[2, 56, 19, 31],\n[41, 18, 6, 45]]");
		$display("Expect: 159, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 38;
		pixel_array_in[0][1] = 60;
		pixel_array_in[0][2] = 8;
		pixel_array_in[0][3] = 43;
		pixel_array_in[1][0] = 19;
		pixel_array_in[1][1] = 11;
		pixel_array_in[1][2] = 4;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 49;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 56;
		pixel_array_in[3][0] = 49;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 1;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[27, 26, 14, 61],\n[47, 6, 49, 45],\n[10, 27, 2, 41],\n[42, 60, 22, 42]]");
		$display("Expect: 32, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 11;
		pixel_array_in[0][2] = 6;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 60;
		pixel_array_in[1][1] = 30;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 11;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 24;
		pixel_array_in[2][2] = 40;
		pixel_array_in[2][3] = 41;
		pixel_array_in[3][0] = 53;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 54;
		#10;
		
		$display("Input: \n[[30, 25, 39, 36],\n[29, 11, 50, 57],\n[42, 53, 58, 42],\n[27, 22, 51, 23]]");
		$display("Expect: 77, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 12;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 25;
		pixel_array_in[1][1] = 16;
		pixel_array_in[1][2] = 23;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 21;
		pixel_array_in[2][1] = 41;
		pixel_array_in[2][2] = 18;
		pixel_array_in[2][3] = 26;
		pixel_array_in[3][0] = 20;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 46;
		pixel_array_in[3][3] = 55;
		#10;
		
		$display("Input: \n[[38, 60, 8, 43],\n[19, 11, 4, 15],\n[49, 10, 22, 56],\n[49, 38, 1, 6]]");
		$display("Expect: 26, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 5;
		pixel_array_in[0][1] = 14;
		pixel_array_in[0][2] = 6;
		pixel_array_in[0][3] = 20;
		pixel_array_in[1][0] = 55;
		pixel_array_in[1][1] = 20;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 14;
		pixel_array_in[2][0] = 54;
		pixel_array_in[2][1] = 40;
		pixel_array_in[2][2] = 41;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 9;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 21;
		#10;
		
		$display("Input: \n[[15, 11, 6, 42],\n[60, 30, 39, 11],\n[47, 24, 40, 41],\n[53, 25, 36, 54]]");
		$display("Expect: 120, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 45;
		pixel_array_in[0][1] = 29;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 7;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 26;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 31;
		pixel_array_in[2][2] = 9;
		pixel_array_in[2][3] = 29;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 2;
		pixel_array_in[3][2] = 25;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[12, 58, 13, 18],\n[25, 16, 23, 48],\n[21, 41, 18, 26],\n[20, 13, 46, 55]]");
		$display("Expect: 75, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 26;
		pixel_array_in[0][1] = 3;
		pixel_array_in[0][2] = 16;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 56;
		pixel_array_in[1][1] = 6;
		pixel_array_in[1][2] = 54;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 23;
		pixel_array_in[2][1] = 52;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 14;
		#10;
		
		$display("Input: \n[[5, 14, 6, 20],\n[55, 20, 25, 14],\n[54, 40, 41, 36],\n[23, 9, 6, 21]]");
		$display("Expect: 100, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 20;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 34;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 22;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 47;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 2;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 52;
		pixel_array_in[3][3] = 53;
		#10;
		
		$display("Input: \n[[45, 29, 55, 7],\n[47, 26, 25, 44],\n[43, 31, 9, 29],\n[29, 2, 25, 39]]");
		$display("Expect: 109, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 43;
		pixel_array_in[0][1] = 16;
		pixel_array_in[0][2] = 29;
		pixel_array_in[0][3] = 53;
		pixel_array_in[1][0] = 26;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 12;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 46;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 29;
		pixel_array_in[2][3] = 34;
		pixel_array_in[3][0] = 4;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[26, 3, 16, 2],\n[56, 6, 54, 17],\n[23, 52, 23, 3],\n[36, 50, 45, 14]]");
		$display("Expect: 62, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 30;
		pixel_array_in[0][1] = 35;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 56;
		pixel_array_in[1][2] = 27;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 28;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 46;
		pixel_array_in[3][0] = 27;
		pixel_array_in[3][1] = 10;
		pixel_array_in[3][2] = 53;
		pixel_array_in[3][3] = 32;
		#10;
		
		$display("Input: \n[[21, 52, 20, 58],\n[58, 34, 32, 22],\n[14, 47, 52, 18],\n[2, 37, 52, 53]]");
		$display("Expect: 142, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 47;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 60;
		pixel_array_in[1][0] = 37;
		pixel_array_in[1][1] = 47;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 43;
		pixel_array_in[2][0] = 25;
		pixel_array_in[2][1] = 21;
		pixel_array_in[2][2] = 3;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 49;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 53;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[43, 16, 29, 53],\n[26, 50, 12, 48],\n[46, 38, 29, 34],\n[4, 48, 51, 44]]");
		$display("Expect: 198, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 52;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 49;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 23;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 24;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 56;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[30, 35, 30, 45],\n[0, 56, 27, 47],\n[28, 3, 17, 46],\n[27, 10, 53, 32]]");
		$display("Expect: 186, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 14;
		pixel_array_in[0][1] = 41;
		pixel_array_in[0][2] = 38;
		pixel_array_in[0][3] = 11;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 61;
		pixel_array_in[1][2] = 51;
		pixel_array_in[1][3] = 50;
		pixel_array_in[2][0] = 19;
		pixel_array_in[2][1] = 26;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 27;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 31;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 15;
		#10;
		
		$display("Input: \n[[19, 47, 12, 60],\n[37, 47, 3, 43],\n[25, 21, 3, 42],\n[49, 28, 53, 1]]");
		$display("Expect: 166, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 18;
		pixel_array_in[0][3] = 35;
		pixel_array_in[1][0] = 33;
		pixel_array_in[1][1] = 15;
		pixel_array_in[1][2] = 59;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 39;
		pixel_array_in[2][2] = 59;
		pixel_array_in[2][3] = 34;
		pixel_array_in[3][0] = 27;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 40;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[52, 7, 49, 41],\n[23, 28, 13, 24],\n[14, 55, 5, 56],\n[15, 37, 2, 7]]");
		$display("Expect: 141, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 41;
		pixel_array_in[0][1] = 14;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 56;
		pixel_array_in[1][0] = 33;
		pixel_array_in[1][1] = 5;
		pixel_array_in[1][2] = 55;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 50;
		pixel_array_in[2][2] = 34;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 8;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[14, 41, 38, 11],\n[11, 61, 51, 50],\n[19, 26, 49, 27],\n[19, 31, 27, 15]]");
		$display("Expect: 220, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 33;
		pixel_array_in[0][1] = 41;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 34;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 5;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 15;
		pixel_array_in[3][2] = 41;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[8, 56, 18, 35],\n[33, 15, 59, 39],\n[39, 39, 59, 34],\n[27, 37, 40, 2]]");
		$display("Expect: 68, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 2;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 20;
		pixel_array_in[0][3] = 26;
		pixel_array_in[1][0] = 8;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 1;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 37;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 7;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 21;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[41, 14, 19, 56],\n[33, 5, 55, 0],\n[24, 50, 34, 18],\n[8, 57, 17, 33]]");
		$display("Expect: 53, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 2;
		pixel_array_in[0][1] = 16;
		pixel_array_in[0][2] = 56;
		pixel_array_in[0][3] = 6;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 16;
		pixel_array_in[1][3] = 1;
		pixel_array_in[2][0] = 59;
		pixel_array_in[2][1] = 27;
		pixel_array_in[2][2] = 16;
		pixel_array_in[2][3] = 12;
		pixel_array_in[3][0] = 8;
		pixel_array_in[3][1] = 1;
		pixel_array_in[3][2] = 58;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[33, 41, 23, 57],\n[34, 54, 37, 15],\n[60, 5, 62, 24],\n[61, 15, 41, 39]]");
		$display("Expect: 178, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 16;
		pixel_array_in[0][1] = 17;
		pixel_array_in[0][2] = 2;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 51;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 25;
		pixel_array_in[2][3] = 33;
		pixel_array_in[3][0] = 11;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 24;
		pixel_array_in[3][3] = 61;
		#10;
		
		$display("Input: \n[[2, 7, 20, 26],\n[8, 50, 37, 1],\n[31, 37, 7, 7],\n[61, 57, 21, 27]]");
		$display("Expect: 199, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 41;
		pixel_array_in[0][3] = 26;
		pixel_array_in[1][0] = 48;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 46;
		pixel_array_in[1][3] = 26;
		pixel_array_in[2][0] = 25;
		pixel_array_in[2][1] = 18;
		pixel_array_in[2][2] = 56;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 28;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 45;
		#10;
		
		$display("Input: \n[[2, 16, 56, 6],\n[44, 32, 16, 1],\n[59, 27, 16, 12],\n[8, 1, 58, 56]]");
		$display("Expect: 130, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 17;
		pixel_array_in[0][1] = 57;
		pixel_array_in[0][2] = 20;
		pixel_array_in[0][3] = 9;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 5;
		pixel_array_in[1][2] = 20;
		pixel_array_in[1][3] = 21;
		pixel_array_in[2][0] = 48;
		pixel_array_in[2][1] = 50;
		pixel_array_in[2][2] = 32;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 50;
		pixel_array_in[3][1] = 29;
		pixel_array_in[3][2] = 44;
		pixel_array_in[3][3] = 30;
		#10;
		
		$display("Input: \n[[16, 17, 2, 36],\n[61, 50, 22, 51],\n[22, 23, 25, 33],\n[11, 42, 24, 61]]");
		$display("Expect: 185, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 5;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 49;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 21;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 34;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 49;
		pixel_array_in[2][2] = 9;
		pixel_array_in[2][3] = 50;
		pixel_array_in[3][0] = 35;
		pixel_array_in[3][1] = 60;
		pixel_array_in[3][2] = 53;
		pixel_array_in[3][3] = 13;
		#10;
		
		$display("Input: \n[[32, 58, 41, 26],\n[48, 23, 46, 26],\n[25, 18, 56, 39],\n[28, 25, 3, 45]]");
		$display("Expect: 77, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 39;
		pixel_array_in[0][1] = 33;
		pixel_array_in[0][2] = 28;
		pixel_array_in[0][3] = 17;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 22;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 31;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 30;
		pixel_array_in[3][1] = 8;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 40;
		#10;
		
		$display("Input: \n[[17, 57, 20, 9],\n[44, 5, 20, 21],\n[48, 50, 32, 55],\n[50, 29, 44, 30]]");
		$display("Expect: 43, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 41;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 57;
		pixel_array_in[1][1] = 55;
		pixel_array_in[1][2] = 9;
		pixel_array_in[1][3] = 5;
		pixel_array_in[2][0] = 58;
		pixel_array_in[2][1] = 8;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 35;
		pixel_array_in[3][0] = 27;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 29;
		#10;
		
		$display("Input: \n[[22, 5, 4, 49],\n[38, 21, 32, 34],\n[43, 49, 9, 50],\n[35, 60, 53, 13]]");
		$display("Expect: 110, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 17;
		pixel_array_in[0][1] = 34;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 13;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 43;
		pixel_array_in[1][2] = 61;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 30;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 50;
		pixel_array_in[3][0] = 22;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[39, 33, 28, 17],\n[9, 22, 5, 47],\n[31, 10, 31, 10],\n[30, 8, 15, 40]]");
		$display("Expect: 75, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 35;
		pixel_array_in[1][1] = 10;
		pixel_array_in[1][2] = 35;
		pixel_array_in[1][3] = 19;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 30;
		pixel_array_in[2][2] = 62;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 56;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 54;
		pixel_array_in[3][3] = 9;
		#10;
		
		$display("Input: \n[[41, 26, 45, 15],\n[57, 55, 9, 5],\n[58, 8, 61, 35],\n[27, 30, 7, 29]]");
		$display("Expect: 187, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 61;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 9;
		pixel_array_in[1][0] = 50;
		pixel_array_in[1][1] = 22;
		pixel_array_in[1][2] = 38;
		pixel_array_in[1][3] = 40;
		pixel_array_in[2][0] = 17;
		pixel_array_in[2][1] = 16;
		pixel_array_in[2][2] = 14;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 35;
		pixel_array_in[3][1] = 35;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 12;
		#10;
		
		$display("Input: \n[[17, 34, 14, 13],\n[32, 43, 61, 48],\n[60, 30, 54, 50],\n[22, 45, 60, 20]]");
		$display("Expect: 162, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 10;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 26;
		pixel_array_in[1][1] = 46;
		pixel_array_in[1][2] = 2;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 37;
		pixel_array_in[3][0] = 62;
		pixel_array_in[3][1] = 60;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 41;
		#10;
		
		$display("Input: \n[[29, 18, 13, 8],\n[35, 10, 35, 19],\n[5, 30, 62, 0],\n[56, 14, 54, 9]]");
		$display("Expect: 55, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 41;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 27;
		pixel_array_in[0][3] = 6;
		pixel_array_in[1][0] = 6;
		pixel_array_in[1][1] = 6;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 33;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 6;
		pixel_array_in[2][2] = 35;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 44;
		pixel_array_in[3][1] = 9;
		pixel_array_in[3][2] = 49;
		pixel_array_in[3][3] = 50;
		#10;
		
		$display("Input: \n[[57, 61, 13, 9],\n[50, 22, 38, 40],\n[17, 16, 14, 62],\n[35, 35, 11, 12]]");
		$display("Expect: 70, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 41;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 59;
		pixel_array_in[0][3] = 34;
		pixel_array_in[1][0] = 3;
		pixel_array_in[1][1] = 22;
		pixel_array_in[1][2] = 40;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 32;
		pixel_array_in[2][1] = 59;
		pixel_array_in[2][2] = 35;
		pixel_array_in[2][3] = 20;
		pixel_array_in[3][0] = 14;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 22;
		pixel_array_in[3][3] = 38;
		#10;
		
		$display("Input: \n[[53, 54, 10, 45],\n[26, 46, 2, 46],\n[39, 1, 5, 37],\n[62, 60, 51, 41]]");
		$display("Expect: 139, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 47;
		pixel_array_in[0][1] = 29;
		pixel_array_in[0][2] = 22;
		pixel_array_in[0][3] = 50;
		pixel_array_in[1][0] = 53;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 16;
		pixel_array_in[1][3] = 11;
		pixel_array_in[2][0] = 51;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 27;
		pixel_array_in[2][3] = 59;
		pixel_array_in[3][0] = 45;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 19;
		#10;
		
		$display("Input: \n[[41, 10, 27, 6],\n[6, 6, 0, 33],\n[40, 6, 35, 24],\n[44, 9, 49, 50]]");
		$display("Expect: 22, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 21;
		pixel_array_in[0][2] = 42;
		pixel_array_in[0][3] = 24;
		pixel_array_in[1][0] = 18;
		pixel_array_in[1][1] = 2;
		pixel_array_in[1][2] = 62;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 26;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 53;
		pixel_array_in[2][3] = 20;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 46;
		pixel_array_in[3][2] = 10;
		pixel_array_in[3][3] = 13;
		#10;
		
		$display("Input: \n[[41, 28, 59, 34],\n[3, 22, 40, 0],\n[32, 59, 35, 20],\n[14, 48, 22, 38]]");
		$display("Expect: 117, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 46;
		pixel_array_in[0][3] = 50;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 24;
		pixel_array_in[1][2] = 9;
		pixel_array_in[1][3] = 8;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 51;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 56;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[47, 29, 22, 50],\n[53, 54, 16, 11],\n[51, 35, 27, 59],\n[45, 25, 3, 19]]");
		$display("Expect: 208, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 51;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 37;
		pixel_array_in[0][3] = 46;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 15;
		pixel_array_in[1][2] = 62;
		pixel_array_in[1][3] = 54;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 34;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 49;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 20;
		#10;
		
		$display("Input: \n[[32, 21, 42, 24],\n[18, 2, 62, 29],\n[26, 10, 53, 20],\n[31, 46, 10, 13]]");
		$display("Expect: 5, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 48;
		pixel_array_in[0][1] = 38;
		pixel_array_in[0][2] = 37;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 19;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 54;
		pixel_array_in[1][3] = 21;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 56;
		pixel_array_in[3][2] = 47;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[29, 45, 46, 50],\n[0, 24, 9, 8],\n[11, 51, 22, 3],\n[23, 56, 32, 7]]");
		$display("Expect: 111, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 7;
		pixel_array_in[0][1] = 62;
		pixel_array_in[0][2] = 35;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 31;
		pixel_array_in[2][1] = 60;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 53;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 46;
		#10;
		
		$display("Input: \n[[51, 28, 37, 46],\n[11, 15, 62, 54],\n[10, 11, 34, 18],\n[49, 34, 27, 20]]");
		$display("Expect: 50, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 46;
		pixel_array_in[0][1] = 45;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 19;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 5;
		pixel_array_in[1][3] = 13;
		pixel_array_in[2][0] = 38;
		pixel_array_in[2][1] = 22;
		pixel_array_in[2][2] = 59;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 2;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 4;
		#10;
		
		$display("Input: \n[[48, 38, 37, 19],\n[19, 35, 54, 21],\n[0, 1, 43, 42],\n[15, 56, 47, 56]]");
		$display("Expect: 106, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 46;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 50;
		pixel_array_in[1][0] = 1;
		pixel_array_in[1][1] = 6;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 52;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 34;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 51;
		#10;
		
		$display("Input: \n[[7, 62, 35, 18],\n[11, 45, 25, 15],\n[31, 60, 52, 62],\n[53, 58, 3, 46]]");
		$display("Expect: 187, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 34;
		pixel_array_in[0][1] = 50;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 37;
		pixel_array_in[1][0] = 2;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 9;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 59;
		pixel_array_in[2][1] = 20;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 26;
		pixel_array_in[3][3] = 57;
		#10;
		
		$display("Input: \n[[46, 45, 4, 58],\n[19, 45, 5, 13],\n[38, 22, 59, 0],\n[29, 2, 56, 4]]");
		$display("Expect: 163, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 59;
		pixel_array_in[0][2] = 44;
		pixel_array_in[0][3] = 11;
		pixel_array_in[1][0] = 34;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 49;
		pixel_array_in[2][0] = 38;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 46;
		pixel_array_in[3][0] = 23;
		pixel_array_in[3][1] = 53;
		pixel_array_in[3][2] = 52;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[46, 54, 14, 50],\n[1, 6, 3, 52],\n[0, 11, 49, 34],\n[52, 6, 59, 51]]");
		$display("Expect: 15, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 18;
		pixel_array_in[0][1] = 61;
		pixel_array_in[0][2] = 2;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 14;
		pixel_array_in[1][1] = 29;
		pixel_array_in[1][2] = 9;
		pixel_array_in[1][3] = 59;
		pixel_array_in[2][0] = 5;
		pixel_array_in[2][1] = 11;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 37;
		pixel_array_in[3][1] = 3;
		pixel_array_in[3][2] = 4;
		pixel_array_in[3][3] = 41;
		#10;
		
		$display("Input: \n[[34, 50, 12, 37],\n[2, 27, 9, 29],\n[59, 20, 19, 49],\n[52, 57, 26, 57]]");
		$display("Expect: 92, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[29, 59, 44, 11],\n[34, 12, 32, 49],\n[38, 13, 49, 46],\n[23, 53, 52, 7]]");
		$display("Expect: 31, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[18, 61, 2, 0],\n[14, 29, 9, 59],\n[5, 11, 7, 44],\n[37, 3, 4, 41]]");
		$display("Expect: 93, Result: %d", pixel_out);
		$display("");
		#10;
		
		
		$display("Finishing Sim"); //print nice message
		$finish;
		
    end
endmodule //counter_tb

`default_nettype wire