`timescale 1ns / 1ps
`default_nettype none

module bicubic_interpolation_tb;
    //make logics for inputs and outputs!
    logic clk_in;
    logic rst_in;
    logic valid_in;
    logic [15:0] pixel_array_in [3:0][3:0];
    logic [7:0] r_out [3:0][3:0];
	logic [7:0] g_out [3:0][3:0];
	logic [7:0] b_out [3:0][3:0];
	logic valid_out;

    bicubic_interpolation uut (
        .clk_in(clk_in),
        .rst_in(rst_in),
		.valid_in(valid_in),
        .pixel_array_in(pixel_array_in),
		.r_out(r_out),
		.g_out(g_out),
		.b_out(b_out),
		.valid_out(valid_out)
    );
    always begin
        #5;  //every 5 ns switch...so period of clock is 10 ns...100 MHz clock
        clk_in = !clk_in;
    end

    //initial block...this is our test simulation
    initial begin
		
		$dumpfile("test/bicubic_interpolation.vcd"); //file to store value change dump (vcd)
		$dumpvars(0,bicubic_interpolation_tb); //store everything at the current level and below
		$display("Starting Sim"); //print nice message
		clk_in = 0; //initialize clk (super important)
		rst_in = 0; //initialize rst (super important)
		
		#10;  //wait a little bit of time at beginning
		rst_in = 1; //reset system
		#10; //hold high for a few clock cycles
		rst_in=0;
		
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 0;
		#10;
		
		pixel_array_in[0][0] = 65535;
		pixel_array_in[0][1] = 65535;
		pixel_array_in[0][2] = 65535;
		pixel_array_in[0][3] = 65535;
		pixel_array_in[1][0] = 65535;
		pixel_array_in[1][1] = 65535;
		pixel_array_in[1][2] = 65535;
		pixel_array_in[1][3] = 65535;
		pixel_array_in[2][0] = 65535;
		pixel_array_in[2][1] = 65535;
		pixel_array_in[2][2] = 65535;
		pixel_array_in[2][3] = 65535;
		pixel_array_in[3][0] = 65535;
		pixel_array_in[3][1] = 65535;
		pixel_array_in[3][2] = 65535;
		pixel_array_in[3][3] = 65535;
		#10;
		
		pixel_array_in[0][0] = 64511;
		pixel_array_in[0][1] = 64511;
		pixel_array_in[0][2] = 64511;
		pixel_array_in[0][3] = 64511;
		pixel_array_in[1][0] = 64511;
		pixel_array_in[1][1] = 64511;
		pixel_array_in[1][2] = 64511;
		pixel_array_in[1][3] = 64511;
		pixel_array_in[2][0] = 64511;
		pixel_array_in[2][1] = 64511;
		pixel_array_in[2][2] = 64511;
		pixel_array_in[2][3] = 64511;
		pixel_array_in[3][0] = 64511;
		pixel_array_in[3][1] = 64511;
		pixel_array_in[3][2] = 64511;
		pixel_array_in[3][3] = 64511;
		#10;
		
		pixel_array_in[0][0] = 65535;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 65535;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 65535;
		pixel_array_in[1][2] = 65535;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 65535;
		pixel_array_in[2][2] = 65535;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 65535;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 65535;
		#10;
		
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 65535;
		pixel_array_in[0][2] = 65535;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 65535;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 65535;
		pixel_array_in[2][0] = 65535;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 65535;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 65535;
		pixel_array_in[3][2] = 65535;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Case 6:");
		$display("\tExpect: \n\t[[0, 0, 0, 0],\t[[0, 0, 0, 0],\t[[0, 0, 0, 0],\n\t[0, 0, 0, 0],\t[0, 0, 0, 0],\t[0, 0, 0, 0],\n\t[0, 0, 0, 0],\t[0, 0, 0, 0],\t[0, 0, 0, 0],\n\t[0, 0, 0, 0]]\t[0, 0, 0, 0]]\t[0, 0, 0, 0]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 61660;
		pixel_array_in[0][1] = 43795;
		pixel_array_in[0][2] = 60897;
		pixel_array_in[0][3] = 15030;
		pixel_array_in[1][0] = 14008;
		pixel_array_in[1][1] = 40525;
		pixel_array_in[1][2] = 13264;
		pixel_array_in[1][3] = 3653;
		pixel_array_in[2][0] = 27133;
		pixel_array_in[2][1] = 44684;
		pixel_array_in[2][2] = 42267;
		pixel_array_in[2][3] = 59511;
		pixel_array_in[3][0] = 57596;
		pixel_array_in[3][1] = 33800;
		pixel_array_in[3][2] = 63329;
		pixel_array_in[3][3] = 24026;
		#10;
		
		$display("Case 7:");
		$display("\tExpect: \n\t[[248, 248, 248, 248],\t[[252, 252, 252, 252],\t[[248, 248, 248, 248],\n\t[248, 248, 248, 248],\t[252, 252, 252, 252],\t[248, 248, 248, 248],\n\t[248, 248, 248, 248],\t[252, 252, 252, 252],\t[248, 248, 248, 248],\n\t[248, 248, 248, 248]]\t[252, 252, 252, 252]]\t[248, 248, 248, 248]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 53043;
		pixel_array_in[0][1] = 41999;
		pixel_array_in[0][2] = 43788;
		pixel_array_in[0][3] = 14372;
		pixel_array_in[1][0] = 23107;
		pixel_array_in[1][1] = 34973;
		pixel_array_in[1][2] = 23949;
		pixel_array_in[1][3] = 59990;
		pixel_array_in[2][0] = 9594;
		pixel_array_in[2][1] = 16592;
		pixel_array_in[2][2] = 17426;
		pixel_array_in[2][3] = 27631;
		pixel_array_in[3][0] = 1999;
		pixel_array_in[3][1] = 10644;
		pixel_array_in[3][2] = 60636;
		pixel_array_in[3][3] = 16465;
		#10;
		
		$display("Case 8:");
		$display("\tExpect: \n\t[[248, 248, 248, 248],\t[[124, 124, 124, 124],\t[[248, 248, 248, 248],\n\t[248, 248, 248, 248],\t[124, 124, 124, 124],\t[248, 248, 248, 248],\n\t[248, 248, 248, 248],\t[124, 124, 124, 124],\t[248, 248, 248, 248],\n\t[248, 248, 248, 248]]\t[124, 124, 124, 124]]\t[248, 248, 248, 248]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 1756;
		pixel_array_in[0][1] = 699;
		pixel_array_in[0][2] = 27863;
		pixel_array_in[0][3] = 931;
		pixel_array_in[1][0] = 60631;
		pixel_array_in[1][1] = 45007;
		pixel_array_in[1][2] = 10876;
		pixel_array_in[1][3] = 37129;
		pixel_array_in[2][0] = 34129;
		pixel_array_in[2][1] = 17877;
		pixel_array_in[2][2] = 58235;
		pixel_array_in[2][3] = 7628;
		pixel_array_in[3][0] = 4865;
		pixel_array_in[3][1] = 12250;
		pixel_array_in[3][2] = 37688;
		pixel_array_in[3][3] = 24035;
		#10;
		
		$display("Case 9:");
		$display("\tExpect: \n\t[[248, 255, 255, 255],\t[[252, 255, 255, 255],\t[[248, 255, 255, 255],\n\t[255, 255, 255, 255],\t[255, 255, 255, 255],\t[255, 255, 255, 255],\n\t[255, 255, 255, 255],\t[255, 255, 255, 255],\t[255, 255, 255, 255],\n\t[255, 255, 255, 255]]\t[255, 255, 255, 255]]\t[255, 255, 255, 255]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 23680;
		pixel_array_in[0][1] = 43411;
		pixel_array_in[0][2] = 17241;
		pixel_array_in[0][3] = 3734;
		pixel_array_in[1][0] = 6373;
		pixel_array_in[1][1] = 15514;
		pixel_array_in[1][2] = 10659;
		pixel_array_in[1][3] = 53292;
		pixel_array_in[2][0] = 36169;
		pixel_array_in[2][1] = 40593;
		pixel_array_in[2][2] = 34012;
		pixel_array_in[2][3] = 52175;
		pixel_array_in[3][0] = 40778;
		pixel_array_in[3][1] = 27206;
		pixel_array_in[3][2] = 58147;
		pixel_array_in[3][3] = 30953;
		#10;
		
		$display("Case 10:");
		$display("\tExpect: \n\t[[0, 0, 0, 0],\t[[0, 0, 0, 0],\t[[0, 0, 0, 0],\n\t[0, 0, 0, 0],\t[0, 0, 0, 0],\t[0, 0, 0, 0],\n\t[0, 0, 0, 0],\t[0, 0, 0, 0],\t[0, 0, 0, 0],\n\t[0, 0, 0, 0]]\t[0, 0, 0, 0]]\t[0, 0, 0, 0]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 51591;
		pixel_array_in[0][1] = 26380;
		pixel_array_in[0][2] = 42572;
		pixel_array_in[0][3] = 33481;
		pixel_array_in[1][0] = 46135;
		pixel_array_in[1][1] = 49393;
		pixel_array_in[1][2] = 7330;
		pixel_array_in[1][3] = 44012;
		pixel_array_in[2][0] = 63240;
		pixel_array_in[2][1] = 2730;
		pixel_array_in[2][2] = 15493;
		pixel_array_in[2][3] = 19372;
		pixel_array_in[3][0] = 59464;
		pixel_array_in[3][1] = 12596;
		pixel_array_in[3][2] = 48778;
		pixel_array_in[3][3] = 18376;
		#10;
		
		$display("Case 11:");
		$display("\tExpect: \n\t[[152, 139, 109, 74],\t[[200, 181, 154, 130],\t[[104, 104, 116, 127],\n\t[155, 142, 112, 78],\t[210, 192, 164, 137],\t[99, 106, 129, 151],\n\t[161, 152, 128, 102],\t[215, 203, 179, 151],\t[99, 112, 144, 177],\n\t[167, 163, 148, 132]]\t[214, 210, 193, 169]]\t[98, 115, 153, 193]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 37548;
		pixel_array_in[0][1] = 59456;
		pixel_array_in[0][2] = 50914;
		pixel_array_in[0][3] = 8206;
		pixel_array_in[1][0] = 10905;
		pixel_array_in[1][1] = 61869;
		pixel_array_in[1][2] = 8547;
		pixel_array_in[1][3] = 30674;
		pixel_array_in[2][0] = 7900;
		pixel_array_in[2][1] = 29078;
		pixel_array_in[2][2] = 42051;
		pixel_array_in[2][3] = 14714;
		pixel_array_in[3][0] = 6731;
		pixel_array_in[3][1] = 33843;
		pixel_array_in[3][2] = 31104;
		pixel_array_in[3][3] = 15770;
		#10;
		
		$display("Case 12:");
		$display("\tExpect: \n\t[[136, 126, 106, 88],\t[[16, 47, 99, 149],\t[[232, 218, 176, 129],\n\t[120, 111, 90, 74],\t[9, 39, 91, 142],\t[218, 206, 170, 131],\n\t[100, 92, 75, 61],\t[11, 34, 80, 127],\t[185, 175, 154, 131],\n\t[79, 75, 64, 55]]\t[18, 34, 71, 111]]\t[149, 143, 138, 133]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 20345;
		pixel_array_in[0][1] = 4456;
		pixel_array_in[0][2] = 1344;
		pixel_array_in[0][3] = 11606;
		pixel_array_in[1][0] = 23114;
		pixel_array_in[1][1] = 19121;
		pixel_array_in[1][2] = 35875;
		pixel_array_in[1][3] = 41654;
		pixel_array_in[2][0] = 36762;
		pixel_array_in[2][1] = 7597;
		pixel_array_in[2][2] = 7782;
		pixel_array_in[2][3] = 12457;
		pixel_array_in[3][0] = 48123;
		pixel_array_in[3][1] = 21527;
		pixel_array_in[3][2] = 56721;
		pixel_array_in[3][3] = 29603;
		#10;
		
		$display("Case 13:");
		$display("\tExpect: \n\t[[168, 135, 93, 57],\t[[248, 220, 170, 116],\t[[120, 140, 177, 212],\n\t[159, 135, 109, 86],\t[245, 218, 168, 114],\t[122, 143, 179, 213],\n\t[128, 125, 128, 133],\t[222, 199, 157, 115],\t[135, 154, 186, 214],\n\t[90, 109, 145, 179]]\t[196, 177, 146, 116]]\t[153, 169, 194, 215]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 52022;
		pixel_array_in[0][1] = 32838;
		pixel_array_in[0][2] = 50166;
		pixel_array_in[0][3] = 22777;
		pixel_array_in[1][0] = 30027;
		pixel_array_in[1][1] = 4292;
		pixel_array_in[1][2] = 15920;
		pixel_array_in[1][3] = 11890;
		pixel_array_in[2][0] = 52421;
		pixel_array_in[2][1] = 43900;
		pixel_array_in[2][2] = 54965;
		pixel_array_in[2][3] = 55187;
		pixel_array_in[3][0] = 42846;
		pixel_array_in[3][1] = 12632;
		pixel_array_in[3][2] = 48711;
		pixel_array_in[3][3] = 3975;
		#10;
		
		$display("Case 14:");
		$display("\tExpect: \n\t[[56, 51, 39, 32],\t[[144, 134, 108, 76],\t[[208, 180, 122, 60],\n\t[68, 63, 52, 45],\t[166, 156, 129, 96],\t[199, 179, 135, 87],\n\t[100, 93, 80, 71],\t[190, 181, 155, 125],\t[181, 178, 162, 140],\n\t[133, 126, 112, 102]]\t[206, 198, 177, 152]]\t[158, 173, 186, 193]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 26048;
		pixel_array_in[0][1] = 10664;
		pixel_array_in[0][2] = 62121;
		pixel_array_in[0][3] = 49443;
		pixel_array_in[1][0] = 63447;
		pixel_array_in[1][1] = 28301;
		pixel_array_in[1][2] = 32981;
		pixel_array_in[1][3] = 40574;
		pixel_array_in[2][0] = 34978;
		pixel_array_in[2][1] = 34099;
		pixel_array_in[2][2] = 7382;
		pixel_array_in[2][3] = 20124;
		pixel_array_in[3][0] = 27269;
		pixel_array_in[3][1] = 27968;
		pixel_array_in[3][2] = 14246;
		pixel_array_in[3][3] = 13309;
		#10;
		
		$display("Case 15:");
		$display("\tExpect: \n\t[[192, 155, 100, 48],\t[[28, 45, 83, 122],\t[[136, 106, 68, 33],\n\t[160, 126, 79, 36],\t[26, 41, 77, 116],\t[125, 98, 61, 30],\n\t[103, 77, 50, 30],\t[46, 55, 84, 118],\t[105, 84, 56, 31],\n\t[44, 29, 26, 30]]\t[71, 75, 97, 124]]\t[86, 73, 54, 36]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 35348;
		pixel_array_in[0][1] = 48412;
		pixel_array_in[0][2] = 62196;
		pixel_array_in[0][3] = 32410;
		pixel_array_in[1][0] = 45260;
		pixel_array_in[1][1] = 51827;
		pixel_array_in[1][2] = 45837;
		pixel_array_in[1][3] = 20530;
		pixel_array_in[2][0] = 18878;
		pixel_array_in[2][1] = 22350;
		pixel_array_in[2][2] = 32964;
		pixel_array_in[2][3] = 31480;
		pixel_array_in[3][0] = 15990;
		pixel_array_in[3][1] = 17622;
		pixel_array_in[3][2] = 22144;
		pixel_array_in[3][3] = 25608;
		#10;
		
		$display("Case 16:");
		$display("\tExpect: \n\t[[240, 209, 143, 73],\t[[52, 43, 33, 30],\t[[104, 78, 50, 29],\n\t[214, 192, 138, 81],\t[52, 44, 38, 38],\t[126, 96, 61, 33],\n\t[175, 168, 141, 109],\t[47, 45, 54, 69],\t[148, 114, 72, 38],\n\t[137, 145, 146, 141]]\t[43, 49, 74, 103]]\t[165, 128, 80, 40]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 10966;
		pixel_array_in[0][1] = 27815;
		pixel_array_in[0][2] = 14743;
		pixel_array_in[0][3] = 40222;
		pixel_array_in[1][0] = 28277;
		pixel_array_in[1][1] = 9181;
		pixel_array_in[1][2] = 38484;
		pixel_array_in[1][3] = 50633;
		pixel_array_in[2][0] = 54685;
		pixel_array_in[2][1] = 15069;
		pixel_array_in[2][2] = 18380;
		pixel_array_in[2][3] = 41007;
		pixel_array_in[3][0] = 40064;
		pixel_array_in[3][1] = 59036;
		pixel_array_in[3][2] = 5966;
		pixel_array_in[3][3] = 54547;
		#10;
		
		$display("Case 17:");
		$display("\tExpect: \n\t[[72, 83, 101, 120],\t[[84, 95, 111, 125],\t[[136, 113, 74, 37],\n\t[64, 72, 87, 104],\t[107, 117, 131, 142],\t[132, 110, 74, 41],\n\t[48, 48, 56, 67],\t[137, 145, 159, 169],\t[119, 98, 68, 42],\n\t[31, 24, 25, 30]]\t[165, 170, 185, 196]]\t[106, 86, 64, 45]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 6949;
		pixel_array_in[0][1] = 54648;
		pixel_array_in[0][2] = 14906;
		pixel_array_in[0][3] = 58037;
		pixel_array_in[1][0] = 52365;
		pixel_array_in[1][1] = 53824;
		pixel_array_in[1][2] = 22670;
		pixel_array_in[1][3] = 5142;
		pixel_array_in[2][0] = 58317;
		pixel_array_in[2][1] = 20033;
		pixel_array_in[2][2] = 61235;
		pixel_array_in[2][3] = 7117;
		pixel_array_in[3][0] = 10072;
		pixel_array_in[3][1] = 3178;
		pixel_array_in[3][2] = 25635;
		pixel_array_in[3][3] = 59566;
		#10;
		
		$display("Case 18:");
		$display("\tExpect: \n\t[[16, 17, 31, 46],\t[[24, 48, 100, 157],\t[[32, 47, 75, 106],\n\t[41, 43, 54, 68],\t[43, 67, 115, 167],\t[70, 83, 102, 121],\n\t[92, 94, 104, 116],\t[71, 92, 133, 177],\t[129, 139, 145, 149],\n\t[142, 146, 156, 167]]\t[96, 114, 148, 185]]\t[186, 193, 187, 174]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 13767;
		pixel_array_in[0][1] = 60990;
		pixel_array_in[0][2] = 57533;
		pixel_array_in[0][3] = 27157;
		pixel_array_in[1][0] = 14820;
		pixel_array_in[1][1] = 15376;
		pixel_array_in[1][2] = 49108;
		pixel_array_in[1][3] = 30477;
		pixel_array_in[2][0] = 46930;
		pixel_array_in[2][1] = 53730;
		pixel_array_in[2][2] = 7055;
		pixel_array_in[2][3] = 43209;
		pixel_array_in[3][0] = 61735;
		pixel_array_in[3][1] = 11977;
		pixel_array_in[3][2] = 35406;
		pixel_array_in[3][3] = 5849;
		#10;
		
		$display("Case 19:");
		$display("\tExpect: \n\t[[104, 98, 106, 118],\t[[208, 163, 102, 47],\t[[104, 109, 126, 148],\n\t[113, 101, 96, 96],\t[209, 172, 115, 65],\t[120, 127, 142, 161],\n\t[121, 104, 86, 73],\t[195, 172, 131, 93],\t[140, 150, 161, 173],\n\t[126, 105, 78, 53]]\t[176, 170, 148, 125]]\t[153, 166, 173, 178]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 20631;
		pixel_array_in[0][1] = 55006;
		pixel_array_in[0][2] = 25324;
		pixel_array_in[0][3] = 46998;
		pixel_array_in[1][0] = 60678;
		pixel_array_in[1][1] = 39133;
		pixel_array_in[1][2] = 29685;
		pixel_array_in[1][3] = 7720;
		pixel_array_in[2][0] = 63188;
		pixel_array_in[2][1] = 28843;
		pixel_array_in[2][2] = 41571;
		pixel_array_in[2][3] = 8375;
		pixel_array_in[3][0] = 34114;
		pixel_array_in[3][1] = 57032;
		pixel_array_in[3][2] = 40683;
		pixel_array_in[3][3] = 941;
		#10;
		
		$display("Case 20:");
		$display("\tExpect: \n\t[[200, 199, 195, 188],\t[[76, 85, 95, 99],\t[[152, 145, 129, 112],\n\t[177, 177, 176, 171],\t[103, 105, 99, 89],\t[137, 126, 108, 92],\n\t[142, 146, 150, 153],\t[153, 141, 110, 74],\t[123, 106, 85, 69],\n\t[105, 114, 124, 134]]\t[203, 178, 122, 62]]\t[113, 90, 65, 48]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 47913;
		pixel_array_in[0][1] = 50336;
		pixel_array_in[0][2] = 30264;
		pixel_array_in[0][3] = 27176;
		pixel_array_in[1][0] = 6035;
		pixel_array_in[1][1] = 60936;
		pixel_array_in[1][2] = 48569;
		pixel_array_in[1][3] = 34098;
		pixel_array_in[2][0] = 8198;
		pixel_array_in[2][1] = 18244;
		pixel_array_in[2][2] = 58988;
		pixel_array_in[2][3] = 27365;
		pixel_array_in[3][0] = 10395;
		pixel_array_in[3][1] = 5979;
		pixel_array_in[3][2] = 47223;
		pixel_array_in[3][3] = 29879;
		#10;
		
		$display("Case 21:");
		$display("\tExpect: \n\t[[32, 48, 80, 116],\t[[120, 130, 155, 182],\t[[232, 223, 205, 182],\n\t[27, 41, 71, 106],\t[108, 126, 163, 201],\t[244, 230, 203, 171],\n\t[29, 34, 58, 88],\t[94, 119, 167, 214],\t[243, 222, 188, 152],\n\t[37, 34, 46, 66]]\t[85, 115, 171, 223]]\t[236, 210, 172, 134]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 40534;
		pixel_array_in[0][1] = 16960;
		pixel_array_in[0][2] = 38149;
		pixel_array_in[0][3] = 34160;
		pixel_array_in[1][0] = 60354;
		pixel_array_in[1][1] = 16097;
		pixel_array_in[1][2] = 16043;
		pixel_array_in[1][3] = 779;
		pixel_array_in[2][0] = 61655;
		pixel_array_in[2][1] = 5289;
		pixel_array_in[2][2] = 10671;
		pixel_array_in[2][3] = 34694;
		pixel_array_in[3][0] = 9758;
		pixel_array_in[3][1] = 23118;
		pixel_array_in[3][2] = 17932;
		pixel_array_in[3][3] = 19913;
		#10;
		
		$display("Case 22:");
		$display("\tExpect: \n\t[[208, 185, 153, 117],\t[[72, 52, 32, 17],\t[[0, 13, 45, 82],\n\t[181, 169, 157, 142],\t[92, 80, 67, 58],\t[0, 3, 41, 84],\n\t[144, 147, 162, 175],\t[133, 131, 128, 126],\t[0, 8, 53, 101],\n\t[104, 121, 163, 202]]\t[175, 184, 190, 192]]\t[0, 21, 69, 119]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 18877;
		pixel_array_in[0][1] = 14837;
		pixel_array_in[0][2] = 51771;
		pixel_array_in[0][3] = 23951;
		pixel_array_in[1][0] = 58752;
		pixel_array_in[1][1] = 178;
		pixel_array_in[1][2] = 49115;
		pixel_array_in[1][3] = 12970;
		pixel_array_in[2][0] = 41841;
		pixel_array_in[2][1] = 29262;
		pixel_array_in[2][2] = 16896;
		pixel_array_in[2][3] = 47458;
		pixel_array_in[3][0] = 25331;
		pixel_array_in[3][1] = 29133;
		pixel_array_in[3][2] = 41615;
		pixel_array_in[3][3] = 8475;
		#10;
		
		$display("Case 23:");
		$display("\tExpect: \n\t[[56, 83, 124, 163],\t[[128, 157, 193, 226],\t[[128, 142, 153, 159],\n\t[78, 92, 113, 133],\t[105, 135, 175, 213],\t[96, 110, 127, 141],\n\t[131, 123, 110, 98],\t[80, 100, 138, 176],\t[61, 75, 100, 124],\n\t[184, 157, 110, 68]]\t[61, 70, 101, 133]]\t[32, 46, 77, 109]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 27543;
		pixel_array_in[0][1] = 32633;
		pixel_array_in[0][2] = 5430;
		pixel_array_in[0][3] = 49076;
		pixel_array_in[1][0] = 52744;
		pixel_array_in[1][1] = 32904;
		pixel_array_in[1][2] = 61713;
		pixel_array_in[1][3] = 44269;
		pixel_array_in[2][0] = 32273;
		pixel_array_in[2][1] = 63145;
		pixel_array_in[2][2] = 1316;
		pixel_array_in[2][3] = 52206;
		pixel_array_in[3][0] = 57276;
		pixel_array_in[3][1] = 748;
		pixel_array_in[3][2] = 36505;
		pixel_array_in[3][3] = 43471;
		#10;
		
		$display("Case 24:");
		$display("\tExpect: \n\t[[152, 140, 132, 124],\t[[24, 33, 61, 95],\t[[232, 234, 218, 192],\n\t[137, 129, 130, 131],\t[5, 13, 45, 84],\t[202, 201, 185, 162],\n\t[122, 118, 128, 139],\t[0, 2, 32, 68],\t[161, 151, 130, 109],\n\t[111, 113, 130, 148]]\t[2, 3, 28, 58]]\t[118, 100, 75, 55]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 37970;
		pixel_array_in[0][1] = 22805;
		pixel_array_in[0][2] = 54539;
		pixel_array_in[0][3] = 41875;
		pixel_array_in[1][0] = 55383;
		pixel_array_in[1][1] = 19978;
		pixel_array_in[1][2] = 2699;
		pixel_array_in[1][3] = 40858;
		pixel_array_in[2][0] = 25031;
		pixel_array_in[2][1] = 7009;
		pixel_array_in[2][2] = 45540;
		pixel_array_in[2][3] = 32924;
		pixel_array_in[3][0] = 41187;
		pixel_array_in[3][1] = 58237;
		pixel_array_in[3][2] = 35448;
		pixel_array_in[3][3] = 45945;
		#10;
		
		$display("Case 25:");
		$display("\tExpect: \n\t[[232, 238, 225, 202],\t[[192, 186, 184, 182],\t[[64, 86, 130, 174],\n\t[201, 216, 216, 208],\t[203, 201, 197, 193],\t[57, 77, 116, 154],\n\t[153, 177, 196, 209],\t[214, 220, 218, 212],\t[40, 58, 91, 124],\n\t[102, 134, 173, 206]]\t[224, 237, 236, 226]]\t[27, 43, 70, 97]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 60985;
		pixel_array_in[0][1] = 63106;
		pixel_array_in[0][2] = 19006;
		pixel_array_in[0][3] = 23427;
		pixel_array_in[1][0] = 57050;
		pixel_array_in[1][1] = 19131;
		pixel_array_in[1][2] = 34557;
		pixel_array_in[1][3] = 5781;
		pixel_array_in[2][0] = 47851;
		pixel_array_in[2][1] = 37637;
		pixel_array_in[2][2] = 11202;
		pixel_array_in[2][3] = 31738;
		pixel_array_in[3][0] = 5467;
		pixel_array_in[3][1] = 48512;
		pixel_array_in[3][2] = 41699;
		pixel_array_in[3][3] = 25469;
		#10;
		
		$display("Case 26:");
		$display("\tExpect: \n\t[[56, 44, 48, 55],\t[[220, 228, 229, 224],\t[[8, 23, 47, 71],\n\t[45, 32, 35, 43],\t[217, 219, 210, 194],\t[20, 35, 59, 83],\n\t[31, 17, 20, 32],\t[198, 192, 168, 141],\t[38, 49, 73, 96],\n\t[18, 4, 10, 25]]\t[171, 158, 123, 88]]\t[56, 63, 84, 106]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 28349;
		pixel_array_in[0][1] = 47896;
		pixel_array_in[0][2] = 60416;
		pixel_array_in[0][3] = 54713;
		pixel_array_in[1][0] = 21164;
		pixel_array_in[1][1] = 39006;
		pixel_array_in[1][2] = 20025;
		pixel_array_in[1][3] = 5873;
		pixel_array_in[2][0] = 44766;
		pixel_array_in[2][1] = 8278;
		pixel_array_in[2][2] = 5122;
		pixel_array_in[2][3] = 40569;
		pixel_array_in[3][0] = 4649;
		pixel_array_in[3][1] = 6343;
		pixel_array_in[3][2] = 55099;
		pixel_array_in[3][3] = 47262;
		#10;
		
		$display("Case 27:");
		$display("\tExpect: \n\t[[0, 24, 86, 150],\t[[20, 59, 134, 209],\t[[144, 171, 197, 214],\n\t[18, 34, 79, 129],\t[28, 61, 126, 190],\t[136, 154, 167, 172],\n\t[52, 54, 74, 99],\t[44, 64, 105, 146],\t[127, 128, 122, 112],\n\t[87, 78, 73, 74]]\t[61, 66, 82, 97]]\t[118, 102, 79, 54]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 28697;
		pixel_array_in[0][1] = 18052;
		pixel_array_in[0][2] = 11218;
		pixel_array_in[0][3] = 10514;
		pixel_array_in[1][0] = 27183;
		pixel_array_in[1][1] = 39258;
		pixel_array_in[1][2] = 56587;
		pixel_array_in[1][3] = 50211;
		pixel_array_in[2][0] = 51430;
		pixel_array_in[2][1] = 26171;
		pixel_array_in[2][2] = 63425;
		pixel_array_in[2][3] = 39128;
		pixel_array_in[3][0] = 15758;
		pixel_array_in[3][1] = 61116;
		pixel_array_in[3][2] = 31219;
		pixel_array_in[3][3] = 5970;
		#10;
		
		$display("Case 28:");
		$display("\tExpect: \n\t[[128, 147, 184, 220],\t[[16, 3, 5, 15],\t[[64, 79, 102, 123],\n\t[156, 164, 180, 195],\t[43, 30, 30, 37],\t[55, 65, 81, 97],\n\t[199, 185, 161, 137],\t[107, 96, 88, 85],\t[58, 57, 60, 65],\n\t[234, 199, 136, 74]]\t[175, 165, 152, 139]]\t[65, 55, 45, 39]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 15921;
		pixel_array_in[0][1] = 13741;
		pixel_array_in[0][2] = 29735;
		pixel_array_in[0][3] = 38578;
		pixel_array_in[1][0] = 15594;
		pixel_array_in[1][1] = 22005;
		pixel_array_in[1][2] = 58823;
		pixel_array_in[1][3] = 36406;
		pixel_array_in[2][0] = 54477;
		pixel_array_in[2][1] = 61644;
		pixel_array_in[2][2] = 53736;
		pixel_array_in[2][3] = 3281;
		pixel_array_in[3][0] = 19665;
		pixel_array_in[3][1] = 45385;
		pixel_array_in[3][2] = 62892;
		pixel_array_in[3][3] = 34720;
		#10;
		
		$display("Case 29:");
		$display("\tExpect: \n\t[[72, 45, 22, 7],\t[[192, 178, 137, 95],\t[[80, 71, 70, 75],\n\t[56, 38, 26, 23],\t[186, 172, 130, 88],\t[53, 46, 47, 56],\n\t[34, 34, 47, 65],\t[160, 148, 116, 81],\t[24, 18, 20, 30],\n\t[19, 37, 74, 113]]\t[128, 120, 100, 77]]\t[4, 0, 1, 11]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 58170;
		pixel_array_in[0][1] = 52100;
		pixel_array_in[0][2] = 26172;
		pixel_array_in[0][3] = 9612;
		pixel_array_in[1][0] = 29694;
		pixel_array_in[1][1] = 20050;
		pixel_array_in[1][2] = 41829;
		pixel_array_in[1][3] = 18644;
		pixel_array_in[2][0] = 62276;
		pixel_array_in[2][1] = 46954;
		pixel_array_in[2][2] = 1993;
		pixel_array_in[2][3] = 59314;
		pixel_array_in[3][0] = 30150;
		pixel_array_in[3][1] = 38100;
		pixel_array_in[3][2] = 33174;
		pixel_array_in[3][3] = 35690;
		#10;
		
		$display("Case 30:");
		$display("\tExpect: \n\t[[72, 75, 98, 121],\t[[84, 102, 144, 190],\t[[216, 221, 228, 233],\n\t[73, 74, 88, 105],\t[75, 95, 137, 181],\t[195, 194, 192, 189],\n\t[95, 84, 81, 81],\t[77, 93, 125, 159],\t[143, 137, 128, 122],\n\t[122, 101, 78, 60]]\t[85, 95, 113, 132]]\t[83, 73, 60, 53]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 5469;
		pixel_array_in[0][1] = 6385;
		pixel_array_in[0][2] = 24099;
		pixel_array_in[0][3] = 30086;
		pixel_array_in[1][0] = 50052;
		pixel_array_in[1][1] = 22890;
		pixel_array_in[1][2] = 21106;
		pixel_array_in[1][3] = 37273;
		pixel_array_in[2][0] = 15752;
		pixel_array_in[2][1] = 8484;
		pixel_array_in[2][2] = 7232;
		pixel_array_in[2][3] = 27574;
		pixel_array_in[3][0] = 13383;
		pixel_array_in[3][1] = 13304;
		pixel_array_in[3][2] = 41463;
		pixel_array_in[3][3] = 26948;
		#10;
		
		$display("Case 31:");
		$display("\tExpect: \n\t[[152, 142, 120, 93],\t[[8, 40, 95, 154],\t[[240, 243, 233, 216],\n\t[125, 111, 88, 63],\t[1, 30, 84, 142],\t[233, 229, 211, 188],\n\t[90, 72, 50, 31],\t[1, 21, 67, 119],\t[218, 198, 162, 127],\n\t[56, 36, 19, 9]]\t[4, 15, 53, 99]]\t[198, 162, 111, 65]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 2829;
		pixel_array_in[0][1] = 42661;
		pixel_array_in[0][2] = 58574;
		pixel_array_in[0][3] = 43300;
		pixel_array_in[1][0] = 30273;
		pixel_array_in[1][1] = 39521;
		pixel_array_in[1][2] = 40526;
		pixel_array_in[1][3] = 42654;
		pixel_array_in[2][0] = 37231;
		pixel_array_in[2][1] = 52497;
		pixel_array_in[2][2] = 29159;
		pixel_array_in[2][3] = 13242;
		pixel_array_in[3][0] = 1626;
		pixel_array_in[3][1] = 38986;
		pixel_array_in[3][2] = 28427;
		pixel_array_in[3][3] = 53287;
		#10;
		
		$display("Case 32:");
		$display("\tExpect: \n\t[[152, 168, 188, 205],\t[[40, 63, 100, 136],\t[[208, 191, 157, 118],\n\t[143, 164, 193, 220],\t[59, 86, 126, 164],\t[221, 198, 151, 100],\n\t[121, 144, 184, 224],\t[106, 136, 175, 207],\t[222, 193, 133, 72],\n\t[99, 125, 172, 221]]\t[159, 190, 223, 245]]\t[217, 184, 116, 48]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 30035;
		pixel_array_in[0][1] = 16193;
		pixel_array_in[0][2] = 56436;
		pixel_array_in[0][3] = 3275;
		pixel_array_in[1][0] = 6491;
		pixel_array_in[1][1] = 16099;
		pixel_array_in[1][2] = 16282;
		pixel_array_in[1][3] = 54752;
		pixel_array_in[2][0] = 45546;
		pixel_array_in[2][1] = 14126;
		pixel_array_in[2][2] = 40982;
		pixel_array_in[2][3] = 935;
		pixel_array_in[3][0] = 6263;
		pixel_array_in[3][1] = 19190;
		pixel_array_in[3][2] = 48171;
		pixel_array_in[3][3] = 35480;
		#10;
		
		$display("Case 33:");
		$display("\tExpect: \n\t[[80, 113, 159, 201],\t[[188, 189, 187, 184],\t[[168, 148, 110, 72],\n\t[116, 143, 181, 214],\t[154, 155, 156, 157],\t[158, 140, 105, 71],\n\t[166, 182, 204, 221],\t[105, 103, 105, 110],\t[137, 122, 94, 67],\n\t[212, 218, 225, 226]]\t[56, 51, 56, 65]]\t[113, 102, 82, 64]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 21385;
		pixel_array_in[0][1] = 2990;
		pixel_array_in[0][2] = 34737;
		pixel_array_in[0][3] = 58407;
		pixel_array_in[1][0] = 57438;
		pixel_array_in[1][1] = 41435;
		pixel_array_in[1][2] = 1676;
		pixel_array_in[1][3] = 48754;
		pixel_array_in[2][0] = 434;
		pixel_array_in[2][1] = 31329;
		pixel_array_in[2][2] = 29775;
		pixel_array_in[2][3] = 46878;
		pixel_array_in[3][0] = 25573;
		pixel_array_in[3][1] = 47298;
		pixel_array_in[3][2] = 23733;
		pixel_array_in[3][3] = 34224;
		#10;
		
		$display("Case 34:");
		$display("\tExpect: \n\t[[72, 89, 119, 147],\t[[200, 188, 164, 134],\t[[144, 113, 78, 50],\n\t[84, 91, 105, 119],\t[215, 207, 185, 158],\t[137, 108, 71, 42],\n\t[118, 103, 88, 77],\t[228, 229, 217, 200],\t[114, 94, 66, 44],\n\t[154, 119, 74, 37]]\t[236, 245, 244, 237]]\t[90, 81, 66, 54]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 37256;
		pixel_array_in[0][1] = 33125;
		pixel_array_in[0][2] = 2445;
		pixel_array_in[0][3] = 22948;
		pixel_array_in[1][0] = 37199;
		pixel_array_in[1][1] = 17904;
		pixel_array_in[1][2] = 9229;
		pixel_array_in[1][3] = 38594;
		pixel_array_in[2][0] = 11174;
		pixel_array_in[2][1] = 12627;
		pixel_array_in[2][2] = 26457;
		pixel_array_in[2][3] = 23696;
		pixel_array_in[3][0] = 3121;
		pixel_array_in[3][1] = 20601;
		pixel_array_in[3][2] = 40651;
		pixel_array_in[3][3] = 50672;
		#10;
		
		$display("Case 35:");
		$display("\tExpect: \n\t[[88, 77, 73, 74],\t[[44, 46, 57, 69],\t[[80, 95, 111, 128],\n\t[80, 68, 62, 61],\t[41, 44, 58, 73],\t[62, 74, 87, 101],\n\t[63, 52, 43, 39],\t[35, 42, 64, 88],\t[42, 44, 47, 53],\n\t[43, 34, 26, 22]]\t[31, 42, 72, 105]]\t[29, 21, 11, 8]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 24616;
		pixel_array_in[0][1] = 59958;
		pixel_array_in[0][2] = 4145;
		pixel_array_in[0][3] = 15750;
		pixel_array_in[1][0] = 42048;
		pixel_array_in[1][1] = 36728;
		pixel_array_in[1][2] = 1006;
		pixel_array_in[1][3] = 55578;
		pixel_array_in[2][0] = 53955;
		pixel_array_in[2][1] = 31636;
		pixel_array_in[2][2] = 18148;
		pixel_array_in[2][3] = 31443;
		pixel_array_in[3][0] = 35846;
		pixel_array_in[3][1] = 35925;
		pixel_array_in[3][2] = 61910;
		pixel_array_in[3][3] = 10821;
		#10;
		
		$display("Case 36:");
		$display("\tExpect: \n\t[[152, 154, 154, 152],\t[[76, 92, 129, 171],\t[[8, 26, 52, 81],\n\t[162, 160, 153, 145],\t[87, 97, 121, 150],\t[33, 43, 57, 75],\n\t[178, 171, 157, 141],\t[119, 118, 117, 118],\t[73, 72, 68, 69],\n\t[193, 182, 162, 139]]\t[150, 140, 115, 89]]\t[113, 101, 80, 64]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 51312;
		pixel_array_in[0][1] = 48576;
		pixel_array_in[0][2] = 37380;
		pixel_array_in[0][3] = 29955;
		pixel_array_in[1][0] = 44448;
		pixel_array_in[1][1] = 135;
		pixel_array_in[1][2] = 34731;
		pixel_array_in[1][3] = 48147;
		pixel_array_in[2][0] = 15484;
		pixel_array_in[2][1] = 47269;
		pixel_array_in[2][2] = 36237;
		pixel_array_in[2][3] = 25044;
		pixel_array_in[3][0] = 204;
		pixel_array_in[3][1] = 20263;
		pixel_array_in[3][2] = 23488;
		pixel_array_in[3][3] = 1780;
		#10;
		
		$display("Case 37:");
		$display("\tExpect: \n\t[[56, 54, 48, 46],\t[[220, 237, 244, 243],\t[[24, 52, 117, 180],\n\t[53, 53, 52, 55],\t[223, 232, 222, 206],\t[41, 69, 127, 183],\n\t[50, 55, 69, 85],\t[231, 220, 184, 142],\t[65, 91, 139, 184],\n\t[47, 59, 90, 120]]\t[235, 206, 144, 79]]\t[90, 112, 149, 180]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 17205;
		pixel_array_in[0][1] = 34870;
		pixel_array_in[0][2] = 63326;
		pixel_array_in[0][3] = 35427;
		pixel_array_in[1][0] = 43383;
		pixel_array_in[1][1] = 30895;
		pixel_array_in[1][2] = 936;
		pixel_array_in[1][3] = 7560;
		pixel_array_in[2][0] = 20852;
		pixel_array_in[2][1] = 17707;
		pixel_array_in[2][2] = 52124;
		pixel_array_in[2][3] = 1900;
		pixel_array_in[3][0] = 23077;
		pixel_array_in[3][1] = 33657;
		pixel_array_in[3][2] = 27419;
		pixel_array_in[3][3] = 4487;
		#10;
		
		$display("Case 38:");
		$display("\tExpect: \n\t[[160, 118, 64, 18],\t[[56, 90, 135, 178],\t[[216, 188, 151, 116],\n\t[161, 125, 75, 32],\t[57, 86, 125, 162],\t[180, 158, 130, 107],\n\t[145, 125, 91, 60],\t[65, 88, 116, 145],\t[118, 106, 98, 96],\n\t[127, 123, 107, 91]]\t[74, 90, 109, 129]]\t[52, 52, 66, 87]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 44360;
		pixel_array_in[0][1] = 53445;
		pixel_array_in[0][2] = 12748;
		pixel_array_in[0][3] = 32209;
		pixel_array_in[1][0] = 33108;
		pixel_array_in[1][1] = 41005;
		pixel_array_in[1][2] = 33549;
		pixel_array_in[1][3] = 51034;
		pixel_array_in[2][0] = 13017;
		pixel_array_in[2][1] = 4449;
		pixel_array_in[2][2] = 39004;
		pixel_array_in[2][3] = 50582;
		pixel_array_in[3][0] = 10313;
		pixel_array_in[3][1] = 62231;
		pixel_array_in[3][2] = 58570;
		pixel_array_in[3][3] = 21035;
		#10;
		
		$display("Case 39:");
		$display("\tExpect: \n\t[[64, 49, 36, 28],\t[[188, 184, 161, 137],\t[[128, 125, 122, 115],\n\t[55, 46, 40, 39],\t[168, 172, 165, 156],\t[137, 139, 139, 135],\n\t[50, 48, 50, 54],\t[124, 140, 158, 174],\t[142, 152, 160, 163],\n\t[47, 52, 61, 71]]\t[75, 103, 146, 189]]\t[145, 162, 177, 187]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 41190;
		pixel_array_in[0][1] = 25029;
		pixel_array_in[0][2] = 13548;
		pixel_array_in[0][3] = 11282;
		pixel_array_in[1][0] = 48728;
		pixel_array_in[1][1] = 37083;
		pixel_array_in[1][2] = 27780;
		pixel_array_in[1][3] = 59459;
		pixel_array_in[2][0] = 4598;
		pixel_array_in[2][1] = 49851;
		pixel_array_in[2][2] = 48168;
		pixel_array_in[2][3] = 17335;
		pixel_array_in[3][0] = 1808;
		pixel_array_in[3][1] = 12996;
		pixel_array_in[3][2] = 6592;
		pixel_array_in[3][3] = 57801;
		#10;
		
		$display("Case 40:");
		$display("\tExpect: \n\t[[136, 101, 53, 11],\t[[236, 222, 192, 155],\t[[192, 187, 158, 126],\n\t[125, 93, 50, 16],\t[222, 217, 201, 180],\t[186, 177, 142, 106],\n\t[121, 91, 55, 27],\t[183, 192, 199, 199],\t[176, 161, 121, 79],\n\t[119, 95, 66, 44]]\t[139, 161, 188, 210]]\t[166, 147, 102, 57]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 3100;
		pixel_array_in[0][1] = 50571;
		pixel_array_in[0][2] = 25184;
		pixel_array_in[0][3] = 62146;
		pixel_array_in[1][0] = 33869;
		pixel_array_in[1][1] = 15220;
		pixel_array_in[1][2] = 24996;
		pixel_array_in[1][3] = 3898;
		pixel_array_in[2][0] = 17322;
		pixel_array_in[2][1] = 49549;
		pixel_array_in[2][2] = 48838;
		pixel_array_in[2][3] = 21344;
		pixel_array_in[3][0] = 10696;
		pixel_array_in[3][1] = 23518;
		pixel_array_in[3][2] = 48688;
		pixel_array_in[3][3] = 17575;
		#10;
		
		$display("Case 41:");
		$display("\tExpect: \n\t[[0, 12, 50, 94],\t[[16, 53, 127, 202],\t[[56, 64, 71, 78],\n\t[27, 39, 68, 103],\t[0, 39, 119, 199],\t[56, 64, 74, 84],\n\t[87, 94, 108, 122],\t[0, 31, 107, 183],\t[50, 55, 70, 89],\n\t[150, 152, 149, 142]]\t[0, 32, 98, 164]]\t[43, 45, 64, 89]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 15692;
		pixel_array_in[0][1] = 51767;
		pixel_array_in[0][2] = 11984;
		pixel_array_in[0][3] = 35405;
		pixel_array_in[1][0] = 1781;
		pixel_array_in[1][1] = 3436;
		pixel_array_in[1][2] = 5174;
		pixel_array_in[1][3] = 54274;
		pixel_array_in[2][0] = 45509;
		pixel_array_in[2][1] = 52010;
		pixel_array_in[2][2] = 36274;
		pixel_array_in[2][3] = 41674;
		pixel_array_in[3][0] = 13907;
		pixel_array_in[3][1] = 54709;
		pixel_array_in[3][2] = 49292;
		pixel_array_in[3][3] = 56436;
		#10;
		
		$display("Case 42:");
		$display("\tExpect: \n\t[[120, 91, 55, 21],\t[[20, 36, 62, 91],\t[[120, 104, 88, 73],\n\t[106, 86, 63, 42],\t[51, 61, 74, 89],\t[106, 97, 91, 88],\n\t[87, 86, 91, 95],\t[96, 100, 98, 98],\t[93, 96, 111, 126],\n\t[70, 90, 123, 152]]\t[139, 137, 123, 110]]\t[85, 102, 137, 171]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 33449;
		pixel_array_in[0][1] = 58205;
		pixel_array_in[0][2] = 30512;
		pixel_array_in[0][3] = 25847;
		pixel_array_in[1][0] = 29396;
		pixel_array_in[1][1] = 24843;
		pixel_array_in[1][2] = 51203;
		pixel_array_in[1][3] = 9589;
		pixel_array_in[2][0] = 57779;
		pixel_array_in[2][1] = 53907;
		pixel_array_in[2][2] = 36089;
		pixel_array_in[2][3] = 10961;
		pixel_array_in[3][0] = 2744;
		pixel_array_in[3][1] = 59909;
		pixel_array_in[3][2] = 23209;
		pixel_array_in[3][3] = 12621;
		#10;
		
		$display("Case 43:");
		$display("\tExpect: \n\t[[160, 154, 142, 130],\t[[4, 16, 39, 66],\t[[104, 97, 94, 95],\n\t[122, 124, 126, 129],\t[9, 17, 31, 52],\t[84, 86, 97, 115],\n\t[71, 82, 100, 121],\t[19, 17, 19, 27],\t[49, 63, 100, 142],\n\t[28, 48, 80, 115]]\t[31, 20, 10, 6]]\t[16, 43, 102, 167]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 48249;
		pixel_array_in[0][1] = 7939;
		pixel_array_in[0][2] = 62281;
		pixel_array_in[0][3] = 43034;
		pixel_array_in[1][0] = 10264;
		pixel_array_in[1][1] = 26187;
		pixel_array_in[1][2] = 5726;
		pixel_array_in[1][3] = 53863;
		pixel_array_in[2][0] = 26443;
		pixel_array_in[2][1] = 62476;
		pixel_array_in[2][2] = 31435;
		pixel_array_in[2][3] = 13147;
		pixel_array_in[3][0] = 9222;
		pixel_array_in[3][1] = 51805;
		pixel_array_in[3][2] = 3852;
		pixel_array_in[3][3] = 42678;
		#10;
		
		$display("Case 44:");
		$display("\tExpect: \n\t[[144, 130, 113, 102],\t[[24, 39, 81, 125],\t[[216, 180, 126, 70],\n\t[160, 153, 139, 129],\t[33, 48, 86, 125],\t[232, 194, 135, 75],\n\t[180, 181, 174, 164],\t[51, 66, 97, 127],\t[238, 201, 142, 83],\n\t[193, 202, 201, 192]]\t[70, 85, 107, 128]]\t[233, 199, 143, 89]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 5747;
		pixel_array_in[0][1] = 25975;
		pixel_array_in[0][2] = 58580;
		pixel_array_in[0][3] = 20824;
		pixel_array_in[1][0] = 44738;
		pixel_array_in[1][1] = 63066;
		pixel_array_in[1][2] = 29451;
		pixel_array_in[1][3] = 938;
		pixel_array_in[2][0] = 48144;
		pixel_array_in[2][1] = 15222;
		pixel_array_in[2][2] = 12387;
		pixel_array_in[2][3] = 29123;
		pixel_array_in[3][0] = 42361;
		pixel_array_in[3][1] = 42383;
		pixel_array_in[3][2] = 42172;
		pixel_array_in[3][3] = 61561;
		#10;
		
		$display("Case 45:");
		$display("\tExpect: \n\t[[56, 61, 77, 92],\t[[108, 90, 67, 50],\t[[160, 133, 88, 46],\n\t[76, 83, 98, 113],\t[89, 82, 75, 75],\t[150, 128, 87, 50],\n\t[122, 129, 138, 144],\t[69, 77, 95, 116],\t[128, 110, 80, 51],\n\t[168, 176, 179, 175]]\t[53, 76, 117, 159]]\t[107, 95, 75, 53]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 32352;
		pixel_array_in[0][1] = 9920;
		pixel_array_in[0][2] = 35816;
		pixel_array_in[0][3] = 44829;
		pixel_array_in[1][0] = 59745;
		pixel_array_in[1][1] = 32398;
		pixel_array_in[1][2] = 21155;
		pixel_array_in[1][3] = 45188;
		pixel_array_in[2][0] = 10466;
		pixel_array_in[2][1] = 56006;
		pixel_array_in[2][2] = 15180;
		pixel_array_in[2][3] = 16744;
		pixel_array_in[3][0] = 27245;
		pixel_array_in[3][1] = 13643;
		pixel_array_in[3][2] = 37253;
		pixel_array_in[3][3] = 53642;
		#10;
		
		$display("Case 46:");
		$display("\tExpect: \n\t[[8, 5, 0, 1],\t[[172, 160, 149, 139],\t[[96, 110, 141, 169],\n\t[33, 30, 24, 24],\t[162, 156, 150, 144],\t[84, 102, 135, 165],\n\t[91, 84, 74, 67],\t[137, 143, 152, 160],\t[77, 96, 128, 156],\n\t[155, 145, 128, 113]]\t[111, 129, 152, 172]]\t[75, 94, 121, 145]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 57769;
		pixel_array_in[0][1] = 48650;
		pixel_array_in[0][2] = 946;
		pixel_array_in[0][3] = 58748;
		pixel_array_in[1][0] = 44778;
		pixel_array_in[1][1] = 57184;
		pixel_array_in[1][2] = 28724;
		pixel_array_in[1][3] = 17222;
		pixel_array_in[2][0] = 38349;
		pixel_array_in[2][1] = 39418;
		pixel_array_in[2][2] = 45481;
		pixel_array_in[2][3] = 18274;
		pixel_array_in[3][0] = 38507;
		pixel_array_in[3][1] = 53520;
		pixel_array_in[3][2] = 2267;
		pixel_array_in[3][3] = 34986;
		#10;
		
		$display("Case 47:");
		$display("\tExpect: \n\t[[96, 119, 157, 190],\t[[32, 17, 1, 0],\t[[88, 66, 42, 25],\n\t[109, 128, 160, 187],\t[37, 26, 15, 10],\t[93, 78, 63, 54],\n\t[142, 150, 166, 178],\t[52, 53, 55, 60],\t[118, 113, 110, 110],\n\t[180, 175, 172, 167]]\t[69, 81, 98, 114]]\t[143, 149, 158, 166]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 20096;
		pixel_array_in[0][1] = 35104;
		pixel_array_in[0][2] = 48140;
		pixel_array_in[0][3] = 1962;
		pixel_array_in[1][0] = 39458;
		pixel_array_in[1][1] = 52626;
		pixel_array_in[1][2] = 13632;
		pixel_array_in[1][3] = 2806;
		pixel_array_in[2][0] = 5178;
		pixel_array_in[2][1] = 43824;
		pixel_array_in[2][2] = 19111;
		pixel_array_in[2][3] = 60177;
		pixel_array_in[3][0] = 15587;
		pixel_array_in[3][1] = 18152;
		pixel_array_in[3][2] = 51505;
		pixel_array_in[3][3] = 49957;
		#10;
		
		$display("Case 48:");
		$display("\tExpect: \n\t[[96, 79, 47, 20],\t[[200, 216, 220, 213],\t[[88, 115, 169, 219],\n\t[131, 112, 73, 36],\t[185, 196, 198, 191],\t[90, 115, 159, 202],\n\t[175, 158, 121, 82],\t[166, 165, 160, 151],\t[87, 102, 130, 158],\n\t[215, 201, 168, 129]]\t[146, 134, 122, 112]]\t[86, 90, 99, 110]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 30482;
		pixel_array_in[0][1] = 30160;
		pixel_array_in[0][2] = 49927;
		pixel_array_in[0][3] = 53602;
		pixel_array_in[1][0] = 26171;
		pixel_array_in[1][1] = 5385;
		pixel_array_in[1][2] = 29990;
		pixel_array_in[1][3] = 18754;
		pixel_array_in[2][0] = 19213;
		pixel_array_in[2][1] = 8090;
		pixel_array_in[2][2] = 52362;
		pixel_array_in[2][3] = 55341;
		pixel_array_in[3][0] = 20932;
		pixel_array_in[3][1] = 24930;
		pixel_array_in[3][2] = 2128;
		pixel_array_in[3][3] = 41455;
		#10;
		
		$display("Case 49:");
		$display("\tExpect: \n\t[[240, 221, 187, 147],\t[[200, 177, 145, 115],\t[[208, 197, 160, 117],\n\t[210, 189, 156, 119],\t[181, 157, 123, 91],\t[204, 188, 146, 98],\n\t[150, 131, 107, 83],\t[151, 126, 92, 60],\t[197, 174, 126, 74],\n\t[89, 74, 61, 54]]\t[122, 98, 65, 34]]\t[187, 159, 109, 56]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 43646;
		pixel_array_in[0][1] = 60260;
		pixel_array_in[0][2] = 18925;
		pixel_array_in[0][3] = 56823;
		pixel_array_in[1][0] = 954;
		pixel_array_in[1][1] = 27652;
		pixel_array_in[1][2] = 32185;
		pixel_array_in[1][3] = 38092;
		pixel_array_in[2][0] = 38653;
		pixel_array_in[2][1] = 40315;
		pixel_array_in[2][2] = 16649;
		pixel_array_in[2][3] = 28793;
		pixel_array_in[3][0] = 58728;
		pixel_array_in[3][1] = 45852;
		pixel_array_in[3][2] = 49596;
		pixel_array_in[3][3] = 54613;
		#10;
		
		$display("Case 50:");
		$display("\tExpect: \n\t[[120, 101, 87, 78],\t[[208, 195, 160, 117],\t[[112, 101, 74, 43],\n\t[149, 127, 101, 78],\t[181, 174, 148, 115],\t[105, 98, 78, 54],\n\t[184, 160, 121, 81],\t[142, 143, 131, 113],\t[84, 85, 79, 69],\n\t[210, 186, 138, 86]]\t[106, 113, 114, 110]]\t[60, 70, 77, 82]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 42769;
		pixel_array_in[0][1] = 10381;
		pixel_array_in[0][2] = 43480;
		pixel_array_in[0][3] = 46255;
		pixel_array_in[1][0] = 4500;
		pixel_array_in[1][1] = 24595;
		pixel_array_in[1][2] = 13463;
		pixel_array_in[1][3] = 46924;
		pixel_array_in[2][0] = 60742;
		pixel_array_in[2][1] = 37877;
		pixel_array_in[2][2] = 28132;
		pixel_array_in[2][3] = 48869;
		pixel_array_in[3][0] = 40121;
		pixel_array_in[3][1] = 56393;
		pixel_array_in[3][2] = 8981;
		pixel_array_in[3][3] = 1422;
		#10;
		
		$display("Case 51:");
		$display("\tExpect: \n\t[[216, 199, 170, 137],\t[[236, 187, 114, 44],\t[[0, 29, 82, 133],\n\t[203, 195, 178, 157],\t[204, 159, 96, 37],\t[38, 58, 93, 126],\n\t[182, 182, 180, 174],\t[152, 118, 74, 36],\t[104, 107, 112, 113],\n\t[161, 168, 178, 182]]\t[98, 76, 52, 37]]\t[169, 157, 133, 104]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 19633;
		pixel_array_in[0][1] = 14097;
		pixel_array_in[0][2] = 5218;
		pixel_array_in[0][3] = 58703;
		pixel_array_in[1][0] = 35843;
		pixel_array_in[1][1] = 35085;
		pixel_array_in[1][2] = 54461;
		pixel_array_in[1][3] = 14524;
		pixel_array_in[2][0] = 48822;
		pixel_array_in[2][1] = 53173;
		pixel_array_in[2][2] = 37377;
		pixel_array_in[2][3] = 29676;
		pixel_array_in[3][0] = 6856;
		pixel_array_in[3][1] = 22300;
		pixel_array_in[3][2] = 54341;
		pixel_array_in[3][3] = 35268;
		#10;
		
		$display("Case 52:");
		$display("\tExpect: \n\t[[200, 173, 129, 82],\t[[176, 183, 183, 177],\t[[144, 119, 69, 19],\n\t[200, 172, 124, 73],\t[167, 173, 171, 164],\t[152, 124, 72, 23],\n\t[194, 169, 120, 70],\t[139, 142, 141, 137],\t[149, 120, 75, 33],\n\t[183, 164, 119, 75]]\t[110, 109, 108, 107]]\t[139, 112, 77, 48]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 22718;
		pixel_array_in[0][1] = 54177;
		pixel_array_in[0][2] = 45482;
		pixel_array_in[0][3] = 58988;
		pixel_array_in[1][0] = 25741;
		pixel_array_in[1][1] = 22162;
		pixel_array_in[1][2] = 32316;
		pixel_array_in[1][3] = 13022;
		pixel_array_in[2][0] = 18607;
		pixel_array_in[2][1] = 54409;
		pixel_array_in[2][2] = 4687;
		pixel_array_in[2][3] = 47474;
		pixel_array_in[3][0] = 11521;
		pixel_array_in[3][1] = 59664;
		pixel_array_in[3][2] = 29170;
		pixel_array_in[3][3] = 11834;
		#10;
		
		$display("Case 53:");
		$display("\tExpect: \n\t[[16, 30, 61, 93],\t[[160, 161, 167, 171],\t[[72, 57, 53, 51],\n\t[9, 28, 66, 105],\t[179, 180, 182, 179],\t[100, 84, 71, 61],\n\t[9, 36, 83, 131],\t[210, 209, 202, 187],\t[148, 129, 103, 77],\n\t[15, 47, 100, 156]]\t[236, 232, 215, 188]]\t[192, 171, 134, 95]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 11268;
		pixel_array_in[0][1] = 17505;
		pixel_array_in[0][2] = 21384;
		pixel_array_in[0][3] = 54341;
		pixel_array_in[1][0] = 57206;
		pixel_array_in[1][1] = 4616;
		pixel_array_in[1][2] = 61116;
		pixel_array_in[1][3] = 38253;
		pixel_array_in[2][0] = 17498;
		pixel_array_in[2][1] = 49039;
		pixel_array_in[2][2] = 29588;
		pixel_array_in[2][3] = 61402;
		pixel_array_in[3][0] = 10627;
		pixel_array_in[3][1] = 55946;
		pixel_array_in[3][2] = 54456;
		pixel_array_in[3][3] = 43914;
		#10;
		
		$display("Case 54:");
		$display("\tExpect: \n\t[[104, 114, 117, 117],\t[[128, 140, 156, 171],\t[[32, 56, 111, 169],\n\t[104, 110, 110, 108],\t[140, 144, 151, 156],\t[69, 82, 117, 156],\n\t[118, 115, 104, 92],\t[156, 147, 135, 123],\t[123, 117, 120, 127],\n\t[137, 124, 101, 79]]\t[168, 145, 116, 86]]\t[178, 153, 124, 100]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 40417;
		pixel_array_in[0][1] = 62165;
		pixel_array_in[0][2] = 4800;
		pixel_array_in[0][3] = 40276;
		pixel_array_in[1][0] = 9990;
		pixel_array_in[1][1] = 6747;
		pixel_array_in[1][2] = 33414;
		pixel_array_in[1][3] = 45539;
		pixel_array_in[2][0] = 41027;
		pixel_array_in[2][1] = 9618;
		pixel_array_in[2][2] = 58702;
		pixel_array_in[2][3] = 53846;
		pixel_array_in[3][0] = 9601;
		pixel_array_in[3][1] = 13364;
		pixel_array_in[3][2] = 28724;
		pixel_array_in[3][3] = 24723;
		#10;
		
		$display("Case 55:");
		$display("\tExpect: \n\t[[96, 88, 69, 50],\t[[0, 23, 63, 107],\t[[152, 160, 173, 183],\n\t[108, 97, 75, 56],\t[23, 47, 85, 126],\t[160, 161, 161, 157],\n\t[119, 106, 88, 74],\t[60, 79, 112, 148],\t[169, 160, 140, 117],\n\t[130, 116, 102, 93]]\t[97, 111, 137, 165]]\t[172, 156, 120, 80]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		pixel_array_in[0][0] = 44591;
		pixel_array_in[0][1] = 49643;
		pixel_array_in[0][2] = 29867;
		pixel_array_in[0][3] = 30361;
		pixel_array_in[1][0] = 20808;
		pixel_array_in[1][1] = 57424;
		pixel_array_in[1][2] = 56403;
		pixel_array_in[1][3] = 58814;
		pixel_array_in[2][0] = 48460;
		pixel_array_in[2][1] = 41381;
		pixel_array_in[2][2] = 10980;
		pixel_array_in[2][3] = 32108;
		pixel_array_in[3][0] = 47981;
		pixel_array_in[3][1] = 51798;
		pixel_array_in[3][2] = 2796;
		pixel_array_in[3][3] = 29163;
		#10;
		
		$display("Case 56:");
		$display("\tExpect: \n\t[[136, 154, 181, 204],\t[[32, 51, 92, 131],\t[[104, 135, 173, 208],\n\t[158, 171, 192, 207],\t[62, 72, 96, 120],\t[113, 136, 160, 184],\n\t[181, 184, 189, 191],\t[127, 119, 113, 108],\t[130, 131, 130, 129],\n\t[197, 191, 181, 169]]\t[197, 172, 134, 98]]\t[150, 129, 98, 70]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		#10;
		
		$display("Case 57:");
		$display("\tExpect: \n\t[[80, 88, 103, 116],\t[[208, 212, 212, 207],\t[[144, 162, 185, 207],\n\t[96, 96, 96, 95],\t[204, 207, 204, 195],\t[137, 155, 176, 196],\n\t[134, 121, 96, 71],\t[188, 189, 178, 161],\t[113, 126, 145, 164],\n\t[177, 151, 101, 52]]\t[167, 164, 146, 121]]\t[85, 93, 111, 129]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		#10;
		
		$display("Case 58:");
		$display("\tExpect: \n\t[[16, 47, 117, 189],\t[[64, 82, 129, 180],\t[[64, 91, 144, 197],\n\t[46, 71, 124, 182],\t[98, 109, 140, 175],\t[80, 102, 149, 196],\n\t[95, 107, 130, 156],\t[157, 154, 155, 159],\t[98, 111, 143, 178],\n\t[146, 144, 137, 131]]\t[213, 197, 169, 142]]\t[112, 117, 135, 158]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		#10;
		
		$display("Case 59:");
		$display("\tExpect: \n\t[[24, 43, 72, 103],\t[[72, 63, 67, 76],\t[[216, 194, 144, 87],\n\t[10, 36, 79, 125],\t[93, 89, 94, 100],\t[204, 187, 144, 97],\n\t[13, 42, 95, 151],\t[125, 130, 135, 137],\t[182, 171, 139, 103],\n\t[24, 54, 112, 173]]\t[157, 168, 172, 169]]\t[158, 154, 132, 109]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		#10;
		
		$display("Case 60:");
		$display("\tExpect: \n\t[[224, 232, 228, 220],\t[[8, 30, 67, 106],\t[[128, 135, 138, 142],\n\t[212, 215, 206, 194],\t[12, 31, 63, 98],\t[109, 115, 117, 121],\n\t[191, 183, 165, 146],\t[25, 36, 60, 89],\t[78, 79, 80, 83],\n\t[170, 151, 122, 94]]\t[40, 43, 59, 80]]\t[49, 45, 44, 46]], \n\tResult:");
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[0][0], r_out[0][1], r_out[0][2], r_out[0][3], g_out[0][0], g_out[0][1], g_out[0][2], g_out[0][3], b_out[0][0], b_out[0][1], b_out[0][2], b_out[0][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[1][0], r_out[1][1], r_out[1][2], r_out[1][3], g_out[1][0], g_out[1][1], g_out[1][2], g_out[1][3], b_out[1][0], b_out[1][1], b_out[1][2], b_out[1][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[2][0], r_out[2][1], r_out[2][2], r_out[2][3], g_out[2][0], g_out[2][1], g_out[2][2], g_out[2][3], b_out[2][0], b_out[2][1], b_out[2][2], b_out[2][3]);
		$display("\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]\t[%d, %d, %d, %d]", r_out[3][0], r_out[3][1], r_out[3][2], r_out[3][3], g_out[3][0], g_out[3][1], g_out[3][2], g_out[3][3], b_out[3][0], b_out[3][1], b_out[3][2], b_out[3][3]);
		$display("");
		#10;
		
		
		$display("Finishing Sim"); //print nice message
		$finish;
		
	end
endmodule //counter_tb

`default_nettype wire