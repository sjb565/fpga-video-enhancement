`timescale 1ns / 1ps
`default_nettype none

module kernel_2_tb;

    //make logics for inputs and outputs!
    logic clk_in;
    logic rst_in;
    logic valid_in;
    logic [5:0] pixel_array_in [3:0][3:0];
    logic [8:0] pixel_out;

    kernel_2 uut (
        .clk_in(clk_in),
        .p1(pixel_array_in[0][1]),
        .p2(pixel_array_in[1][1]),
        .p3(pixel_array_in[2][1]),
        .p4(pixel_array_in[3][1]),
        .pixel_out(pixel_out)
    );
    always begin
        #5;  //every 5 ns switch...so period of clock is 10 ns...100 MHz clock
        clk_in = !clk_in;
    end

    //initial block...this is our test simulation
    initial begin
        
		$dumpfile("test/kernel_2.vcd"); //file to store value change dump (vcd)
		$dumpvars(0,kernel_2_tb); //store everything at the current level and below
		$display("Starting Sim"); //print nice message
		clk_in = 0; //initialize clk (super important)
		rst_in = 0; //initialize rst (super important)
		
		#10;  //wait a little bit of time at beginning
		rst_in = 1; //reset system
		#10; //hold high for a few clock cycles
		rst_in=0;
		
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 0;
		#10;
		
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 32;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 32;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 32;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 32;
		#10;
		
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 63;
		#10;
		
		$display("Input: \n[[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0],\n[0, 0, 0, 0]]");
		$display("Expect: 0, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 63;
		pixel_array_in[0][1] = 0;
		pixel_array_in[0][2] = 0;
		pixel_array_in[0][3] = 63;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 63;
		pixel_array_in[1][2] = 63;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 63;
		pixel_array_in[2][2] = 63;
		pixel_array_in[2][3] = 0;
		pixel_array_in[3][0] = 63;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 0;
		pixel_array_in[3][3] = 63;
		#10;
		
		$display("Input: \n[[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32],\n[32, 32, 32, 32]]");
		$display("Expect: 128, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 63;
		pixel_array_in[0][2] = 63;
		pixel_array_in[0][3] = 0;
		pixel_array_in[1][0] = 63;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 0;
		pixel_array_in[1][3] = 63;
		pixel_array_in[2][0] = 63;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 63;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 63;
		pixel_array_in[3][2] = 63;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Input: \n[[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63],\n[63, 63, 63, 63]]");
		$display("Expect: 252, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 4;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 39;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 55;
		pixel_array_in[1][2] = 28;
		pixel_array_in[1][3] = 55;
		pixel_array_in[2][0] = 13;
		pixel_array_in[2][1] = 9;
		pixel_array_in[2][2] = 29;
		pixel_array_in[2][3] = 20;
		pixel_array_in[3][0] = 9;
		pixel_array_in[3][1] = 59;
		pixel_array_in[3][2] = 62;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[63, 0, 0, 63],\n[0, 63, 63, 0],\n[0, 63, 63, 0],\n[63, 0, 0, 63]]");
		$display("Expect: 384>val>255, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 44;
		pixel_array_in[0][1] = 6;
		pixel_array_in[0][2] = 31;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 36;
		pixel_array_in[1][1] = 8;
		pixel_array_in[1][2] = 27;
		pixel_array_in[1][3] = 58;
		pixel_array_in[2][0] = 24;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 20;
		pixel_array_in[3][3] = 53;
		#10;
		
		$display("Input: \n[[0, 63, 63, 0],\n[63, 0, 0, 63],\n[63, 0, 0, 63],\n[0, 63, 63, 0]]");
		$display("Expect: val>383, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 59;
		pixel_array_in[0][2] = 43;
		pixel_array_in[0][3] = 28;
		pixel_array_in[1][0] = 54;
		pixel_array_in[1][1] = 51;
		pixel_array_in[1][2] = 61;
		pixel_array_in[1][3] = 61;
		pixel_array_in[2][0] = 20;
		pixel_array_in[2][1] = 49;
		pixel_array_in[2][2] = 14;
		pixel_array_in[2][3] = 61;
		pixel_array_in[3][0] = 34;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 12;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[4, 32, 19, 39],\n[0, 55, 28, 55],\n[13, 9, 29, 20],\n[9, 59, 62, 56]]");
		$display("Expect: 121, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 6;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 41;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 23;
		pixel_array_in[1][3] = 14;
		pixel_array_in[2][0] = 51;
		pixel_array_in[2][1] = 26;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 58;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[44, 6, 31, 55],\n[36, 8, 27, 58],\n[24, 10, 5, 42],\n[15, 55, 20, 53]]");
		$display("Expect: 25, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 42;
		pixel_array_in[0][2] = 27;
		pixel_array_in[0][3] = 29;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 18;
		pixel_array_in[1][2] = 24;
		pixel_array_in[1][3] = 50;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 13;
		pixel_array_in[2][3] = 56;
		pixel_array_in[3][0] = 30;
		pixel_array_in[3][1] = 12;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 13;
		#10;
		
		$display("Input: \n[[61, 59, 43, 28],\n[54, 51, 61, 61],\n[20, 49, 14, 61],\n[34, 38, 12, 16]]");
		$display("Expect: 200, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 55;
		pixel_array_in[0][1] = 14;
		pixel_array_in[0][2] = 1;
		pixel_array_in[0][3] = 12;
		pixel_array_in[1][0] = 26;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 11;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 55;
		pixel_array_in[2][1] = 20;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 8;
		pixel_array_in[3][0] = 54;
		pixel_array_in[3][1] = 5;
		pixel_array_in[3][2] = 5;
		pixel_array_in[3][3] = 36;
		#10;
		
		$display("Input: \n[[1, 25, 6, 25],\n[41, 49, 23, 14],\n[51, 26, 42, 36],\n[58, 14, 45, 2]]");
		$display("Expect: 159, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 27;
		pixel_array_in[0][2] = 11;
		pixel_array_in[0][3] = 56;
		pixel_array_in[1][0] = 37;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 61;
		pixel_array_in[1][3] = 41;
		pixel_array_in[2][0] = 8;
		pixel_array_in[2][1] = 58;
		pixel_array_in[2][2] = 53;
		pixel_array_in[2][3] = 13;
		pixel_array_in[3][0] = 57;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 38;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[57, 42, 27, 29],\n[22, 18, 24, 50],\n[50, 1, 13, 56],\n[30, 12, 15, 13]]");
		$display("Expect: 29, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 7;
		pixel_array_in[0][1] = 50;
		pixel_array_in[0][2] = 41;
		pixel_array_in[0][3] = 9;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 38;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 13;
		pixel_array_in[2][1] = 4;
		pixel_array_in[2][2] = 46;
		pixel_array_in[2][3] = 51;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 3;
		pixel_array_in[3][2] = 40;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[55, 14, 1, 12],\n[26, 60, 11, 15],\n[55, 20, 54, 8],\n[54, 5, 5, 36]]");
		$display("Expect: 175, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 35;
		pixel_array_in[0][1] = 51;
		pixel_array_in[0][2] = 52;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 19;
		pixel_array_in[1][3] = 58;
		pixel_array_in[2][0] = 29;
		pixel_array_in[2][1] = 54;
		pixel_array_in[2][2] = 50;
		pixel_array_in[2][3] = 1;
		pixel_array_in[3][0] = 30;
		pixel_array_in[3][1] = 41;
		pixel_array_in[3][2] = 13;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[1, 27, 11, 56],\n[37, 32, 61, 41],\n[8, 58, 53, 13],\n[57, 30, 38, 6]]");
		$display("Expect: 188, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 36;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 48;
		pixel_array_in[1][0] = 15;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 47;
		pixel_array_in[1][3] = 14;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 59;
		pixel_array_in[2][2] = 28;
		pixel_array_in[2][3] = 42;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 57;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[7, 50, 41, 9],\n[44, 38, 36, 15],\n[13, 4, 46, 51],\n[15, 3, 40, 16]]");
		$display("Expect: 81, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 38;
		pixel_array_in[0][1] = 20;
		pixel_array_in[0][2] = 35;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 36;
		pixel_array_in[1][2] = 31;
		pixel_array_in[1][3] = 29;
		pixel_array_in[2][0] = 45;
		pixel_array_in[2][1] = 29;
		pixel_array_in[2][2] = 48;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 26;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 62;
		#10;
		
		$display("Input: \n[[35, 51, 52, 25],\n[28, 28, 19, 58],\n[29, 54, 50, 1],\n[30, 41, 13, 1]]");
		$display("Expect: 161, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 49;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 18;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 46;
		pixel_array_in[1][3] = 42;
		pixel_array_in[2][0] = 62;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 48;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 56;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[9, 36, 14, 48],\n[15, 7, 47, 14],\n[12, 59, 28, 42],\n[42, 57, 36, 27]]");
		$display("Expect: 125, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 41;
		pixel_array_in[0][1] = 21;
		pixel_array_in[0][2] = 14;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 45;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 6;
		pixel_array_in[1][3] = 19;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 0;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 5;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 3;
		pixel_array_in[3][2] = 46;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[38, 20, 35, 25],\n[32, 36, 31, 29],\n[45, 29, 48, 49],\n[26, 25, 15, 62]]");
		$display("Expect: 135, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 54;
		pixel_array_in[0][1] = 39;
		pixel_array_in[0][2] = 29;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 55;
		pixel_array_in[1][2] = 40;
		pixel_array_in[1][3] = 23;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 2;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 45;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 39;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[15, 49, 34, 45],\n[18, 33, 46, 42],\n[62, 12, 48, 18],\n[36, 6, 56, 6]]");
		$display("Expect: 87, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 35;
		pixel_array_in[0][1] = 50;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 51;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 1;
		pixel_array_in[1][3] = 60;
		pixel_array_in[2][0] = 46;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 56;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[41, 21, 14, 36],\n[45, 32, 6, 19],\n[1, 0, 19, 5],\n[42, 3, 46, 39]]");
		$display("Expect: 66, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 37;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 61;
		pixel_array_in[0][3] = 19;
		pixel_array_in[1][0] = 53;
		pixel_array_in[1][1] = 0;
		pixel_array_in[1][2] = 15;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 18;
		pixel_array_in[2][1] = 52;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 55;
		pixel_array_in[3][1] = 5;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 22;
		#10;
		
		$display("Input: \n[[54, 39, 29, 45],\n[31, 55, 40, 23],\n[43, 2, 22, 45],\n[36, 34, 39, 27]]");
		$display("Expect: 110, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 57;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 55;
		pixel_array_in[1][1] = 20;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 28;
		pixel_array_in[2][0] = 4;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 34;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 48;
		pixel_array_in[3][1] = 16;
		pixel_array_in[3][2] = 20;
		pixel_array_in[3][3] = 54;
		#10;
		
		$display("Input: \n[[35, 50, 32, 55],\n[51, 37, 1, 60],\n[46, 10, 23, 3],\n[56, 26, 11, 16]]");
		$display("Expect: 86, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 3;
		pixel_array_in[0][2] = 56;
		pixel_array_in[0][3] = 29;
		pixel_array_in[1][0] = 42;
		pixel_array_in[1][1] = 16;
		pixel_array_in[1][2] = 54;
		pixel_array_in[1][3] = 51;
		pixel_array_in[2][0] = 16;
		pixel_array_in[2][1] = 41;
		pixel_array_in[2][2] = 39;
		pixel_array_in[2][3] = 48;
		pixel_array_in[3][0] = 7;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 21;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[37, 48, 61, 19],\n[53, 0, 15, 15],\n[18, 52, 17, 10],\n[55, 5, 32, 22]]");
		$display("Expect: 103, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 16;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 6;
		pixel_array_in[0][3] = 9;
		pixel_array_in[1][0] = 5;
		pixel_array_in[1][1] = 20;
		pixel_array_in[1][2] = 60;
		pixel_array_in[1][3] = 31;
		pixel_array_in[2][0] = 20;
		pixel_array_in[2][1] = 2;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 54;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 20;
		pixel_array_in[3][2] = 57;
		pixel_array_in[3][3] = 47;
		#10;
		
		$display("Input: \n[[57, 19, 23, 8],\n[55, 20, 39, 28],\n[4, 38, 34, 30],\n[48, 16, 20, 54]]");
		$display("Expect: 121, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 37;
		pixel_array_in[0][2] = 42;
		pixel_array_in[0][3] = 16;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 17;
		pixel_array_in[1][3] = 23;
		pixel_array_in[2][0] = 47;
		pixel_array_in[2][1] = 50;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 2;
		pixel_array_in[3][0] = 22;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 24;
		pixel_array_in[3][3] = 10;
		#10;
		
		$display("Input: \n[[53, 3, 56, 29],\n[42, 16, 54, 51],\n[16, 41, 39, 48],\n[7, 26, 21, 35]]");
		$display("Expect: 121, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 3;
		pixel_array_in[0][2] = 31;
		pixel_array_in[0][3] = 30;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 4;
		pixel_array_in[1][2] = 51;
		pixel_array_in[1][3] = 42;
		pixel_array_in[2][0] = 35;
		pixel_array_in[2][1] = 2;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 58;
		pixel_array_in[3][0] = 3;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 8;
		#10;
		
		$display("Input: \n[[16, 32, 6, 9],\n[5, 20, 60, 31],\n[20, 2, 54, 54],\n[17, 20, 57, 47]]");
		$display("Expect: 36, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 14;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 25;
		pixel_array_in[0][3] = 16;
		pixel_array_in[1][0] = 18;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 44;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 28;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 37;
		pixel_array_in[2][3] = 57;
		pixel_array_in[3][0] = 11;
		pixel_array_in[3][1] = 40;
		pixel_array_in[3][2] = 9;
		pixel_array_in[3][3] = 36;
		#10;
		
		$display("Input: \n[[25, 37, 42, 16],\n[32, 52, 17, 23],\n[47, 50, 49, 2],\n[22, 18, 24, 10]]");
		$display("Expect: 215, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 47;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 57;
		pixel_array_in[0][3] = 4;
		pixel_array_in[1][0] = 40;
		pixel_array_in[1][1] = 41;
		pixel_array_in[1][2] = 28;
		pixel_array_in[1][3] = 42;
		pixel_array_in[2][0] = 19;
		pixel_array_in[2][1] = 16;
		pixel_array_in[2][2] = 10;
		pixel_array_in[2][3] = 11;
		pixel_array_in[3][0] = 9;
		pixel_array_in[3][1] = 11;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 14;
		#10;
		
		$display("Input: \n[[53, 3, 31, 30],\n[13, 4, 51, 42],\n[35, 2, 17, 58],\n[3, 34, 6, 8]]");
		$display("Expect: 4, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 17;
		pixel_array_in[0][1] = 10;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 2;
		pixel_array_in[1][1] = 21;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 54;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 11;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 5;
		pixel_array_in[3][2] = 22;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[14, 19, 25, 16],\n[18, 37, 44, 47],\n[28, 36, 37, 57],\n[11, 40, 9, 36]]");
		$display("Expect: 149, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 46;
		pixel_array_in[0][1] = 35;
		pixel_array_in[0][2] = 58;
		pixel_array_in[0][3] = 7;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 48;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 12;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 51;
		pixel_array_in[2][2] = 12;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 7;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 30;
		pixel_array_in[3][3] = 60;
		#10;
		
		$display("Input: \n[[47, 26, 57, 4],\n[40, 41, 28, 42],\n[19, 16, 10, 11],\n[9, 11, 3, 14]]");
		$display("Expect: 119, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 37;
		pixel_array_in[0][1] = 44;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 18;
		pixel_array_in[1][0] = 45;
		pixel_array_in[1][1] = 6;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 58;
		pixel_array_in[2][1] = 34;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 62;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 2;
		pixel_array_in[3][2] = 20;
		pixel_array_in[3][3] = 0;
		#10;
		
		$display("Input: \n[[17, 10, 30, 45],\n[2, 21, 13, 54],\n[12, 32, 54, 11],\n[61, 5, 22, 52]]");
		$display("Expect: 115, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 16;
		pixel_array_in[0][1] = 27;
		pixel_array_in[0][2] = 5;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 21;
		pixel_array_in[2][0] = 11;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 17;
		pixel_array_in[2][3] = 57;
		pixel_array_in[3][0] = 56;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[46, 35, 58, 7],\n[58, 48, 25, 12],\n[11, 51, 12, 43],\n[7, 25, 30, 60]]");
		$display("Expect: 207, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 56;
		pixel_array_in[0][3] = 10;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 11;
		pixel_array_in[1][2] = 48;
		pixel_array_in[1][3] = 7;
		pixel_array_in[2][0] = 7;
		pixel_array_in[2][1] = 57;
		pixel_array_in[2][2] = 36;
		pixel_array_in[2][3] = 5;
		pixel_array_in[3][0] = 21;
		pixel_array_in[3][1] = 26;
		pixel_array_in[3][2] = 41;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[37, 44, 4, 18],\n[45, 6, 50, 38],\n[58, 34, 17, 62],\n[41, 2, 20, 0]]");
		$display("Expect: 78, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 30;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 34;
		pixel_array_in[1][0] = 2;
		pixel_array_in[1][1] = 28;
		pixel_array_in[1][2] = 53;
		pixel_array_in[1][3] = 51;
		pixel_array_in[2][0] = 3;
		pixel_array_in[2][1] = 1;
		pixel_array_in[2][2] = 28;
		pixel_array_in[2][3] = 10;
		pixel_array_in[3][0] = 26;
		pixel_array_in[3][1] = 39;
		pixel_array_in[3][2] = 54;
		pixel_array_in[3][3] = 59;
		#10;
		
		$display("Input: \n[[16, 27, 5, 36],\n[44, 33, 56, 21],\n[11, 12, 17, 57],\n[56, 58, 11, 1]]");
		$display("Expect: 80, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 29;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 29;
		pixel_array_in[1][0] = 40;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 16;
		pixel_array_in[1][3] = 22;
		pixel_array_in[2][0] = 62;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 29;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 26;
		pixel_array_in[3][3] = 24;
		#10;
		
		$display("Input: \n[[15, 58, 56, 10],\n[31, 11, 48, 7],\n[7, 57, 36, 5],\n[21, 26, 41, 44]]");
		$display("Expect: 132, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 47;
		pixel_array_in[0][1] = 50;
		pixel_array_in[0][2] = 60;
		pixel_array_in[0][3] = 36;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 4;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 13;
		pixel_array_in[2][1] = 42;
		pixel_array_in[2][2] = 12;
		pixel_array_in[2][3] = 17;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 44;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 47;
		#10;
		
		$display("Input: \n[[22, 30, 4, 34],\n[2, 28, 53, 51],\n[3, 1, 28, 10],\n[26, 39, 54, 59]]");
		$display("Expect: 48, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 43;
		pixel_array_in[0][2] = 44;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 14;
		pixel_array_in[1][1] = 43;
		pixel_array_in[1][2] = 57;
		pixel_array_in[1][3] = 8;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 41;
		pixel_array_in[2][2] = 50;
		pixel_array_in[2][3] = 36;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 55;
		pixel_array_in[3][2] = 43;
		pixel_array_in[3][3] = 59;
		#10;
		
		$display("Input: \n[[29, 58, 30, 29],\n[40, 27, 16, 22],\n[62, 3, 29, 44],\n[29, 58, 26, 24]]");
		$display("Expect: 38, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 31;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 57;
		pixel_array_in[0][3] = 30;
		pixel_array_in[1][0] = 26;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 23;
		pixel_array_in[1][3] = 37;
		pixel_array_in[2][0] = 34;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 16;
		pixel_array_in[2][3] = 23;
		pixel_array_in[3][0] = 16;
		pixel_array_in[3][1] = 41;
		pixel_array_in[3][2] = 43;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[47, 50, 60, 36],\n[9, 4, 32, 4],\n[13, 42, 12, 17],\n[52, 44, 60, 47]]");
		$display("Expect: 80, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 20;
		pixel_array_in[0][2] = 1;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 53;
		pixel_array_in[2][0] = 0;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 38;
		pixel_array_in[3][1] = 33;
		pixel_array_in[3][2] = 4;
		pixel_array_in[3][3] = 31;
		#10;
		
		$display("Input: \n[[32, 43, 44, 25],\n[14, 43, 57, 8],\n[14, 41, 50, 36],\n[46, 55, 43, 59]]");
		$display("Expect: 164, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 58;
		pixel_array_in[0][2] = 9;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 21;
		pixel_array_in[1][1] = 44;
		pixel_array_in[1][2] = 60;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 31;
		pixel_array_in[2][2] = 8;
		pixel_array_in[2][3] = 21;
		pixel_array_in[3][0] = 55;
		pixel_array_in[3][1] = 21;
		pixel_array_in[3][2] = 3;
		pixel_array_in[3][3] = 55;
		#10;
		
		$display("Input: \n[[31, 58, 57, 30],\n[26, 35, 23, 37],\n[34, 36, 16, 23],\n[16, 41, 43, 35]]");
		$display("Expect: 135, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 15;
		pixel_array_in[0][3] = 13;
		pixel_array_in[1][0] = 16;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 53;
		pixel_array_in[1][3] = 45;
		pixel_array_in[2][0] = 60;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 30;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 38;
		pixel_array_in[3][3] = 57;
		#10;
		
		$display("Input: \n[[15, 20, 1, 59],\n[9, 35, 3, 53],\n[0, 13, 7, 30],\n[38, 33, 4, 31]]");
		$display("Expect: 94, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 21;
		pixel_array_in[0][2] = 11;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 24;
		pixel_array_in[1][1] = 2;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 57;
		pixel_array_in[2][0] = 39;
		pixel_array_in[2][1] = 55;
		pixel_array_in[2][2] = 29;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 54;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 24;
		#10;
		
		$display("Input: \n[[21, 58, 9, 1],\n[21, 44, 60, 44],\n[12, 31, 8, 21],\n[55, 21, 3, 55]]");
		$display("Expect: 149, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 30;
		pixel_array_in[0][1] = 59;
		pixel_array_in[0][2] = 18;
		pixel_array_in[0][3] = 23;
		pixel_array_in[1][0] = 27;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 26;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 49;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 61;
		pixel_array_in[3][0] = 17;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 14;
		pixel_array_in[3][3] = 38;
		#10;
		
		$display("Input: \n[[61, 52, 15, 13],\n[16, 52, 53, 45],\n[60, 23, 30, 39],\n[36, 18, 38, 57]]");
		$display("Expect: 151, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 44;
		pixel_array_in[0][1] = 6;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 8;
		pixel_array_in[1][1] = 47;
		pixel_array_in[1][2] = 10;
		pixel_array_in[1][3] = 5;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 38;
		pixel_array_in[2][2] = 18;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 3;
		pixel_array_in[3][1] = 51;
		pixel_array_in[3][2] = 14;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[22, 21, 11, 15],\n[24, 2, 22, 57],\n[39, 55, 29, 39],\n[54, 34, 6, 24]]");
		$display("Expect: 114, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 21;
		pixel_array_in[0][3] = 9;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 1;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 4;
		pixel_array_in[2][1] = 36;
		pixel_array_in[2][2] = 10;
		pixel_array_in[2][3] = 54;
		pixel_array_in[3][0] = 41;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 25;
		pixel_array_in[3][3] = 57;
		#10;
		
		$display("Input: \n[[30, 59, 18, 23],\n[27, 50, 26, 4],\n[49, 35, 44, 61],\n[17, 45, 14, 38]]");
		$display("Expect: 165, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 32;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 22;
		pixel_array_in[0][3] = 17;
		pixel_array_in[1][0] = 2;
		pixel_array_in[1][1] = 59;
		pixel_array_in[1][2] = 8;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 33;
		pixel_array_in[2][1] = 37;
		pixel_array_in[2][2] = 11;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 28;
		pixel_array_in[3][1] = 36;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 45;
		#10;
		
		$display("Input: \n[[44, 6, 45, 40],\n[8, 47, 10, 5],\n[15, 38, 18, 18],\n[3, 51, 14, 42]]");
		$display("Expect: 177, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 35;
		pixel_array_in[0][1] = 26;
		pixel_array_in[0][2] = 43;
		pixel_array_in[0][3] = 9;
		pixel_array_in[1][0] = 34;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 44;
		pixel_array_in[1][3] = 39;
		pixel_array_in[2][0] = 54;
		pixel_array_in[2][1] = 58;
		pixel_array_in[2][2] = 58;
		pixel_array_in[2][3] = 58;
		pixel_array_in[3][0] = 21;
		pixel_array_in[3][1] = 5;
		pixel_array_in[3][2] = 53;
		pixel_array_in[3][3] = 17;
		#10;
		
		$display("Input: \n[[19, 18, 21, 9],\n[47, 45, 1, 47],\n[4, 36, 10, 54],\n[41, 0, 25, 57]]");
		$display("Expect: 177, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 5;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 53;
		pixel_array_in[0][3] = 62;
		pixel_array_in[1][0] = 4;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 28;
		pixel_array_in[1][3] = 31;
		pixel_array_in[2][0] = 33;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 33;
		pixel_array_in[2][3] = 60;
		pixel_array_in[3][0] = 21;
		pixel_array_in[3][1] = 23;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 37;
		#10;
		
		$display("Input: \n[[32, 7, 22, 17],\n[2, 59, 8, 47],\n[33, 37, 11, 44],\n[28, 36, 29, 45]]");
		$display("Expect: 205, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 25;
		pixel_array_in[0][1] = 55;
		pixel_array_in[0][2] = 44;
		pixel_array_in[0][3] = 62;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 37;
		pixel_array_in[1][3] = 19;
		pixel_array_in[2][0] = 6;
		pixel_array_in[2][1] = 53;
		pixel_array_in[2][2] = 6;
		pixel_array_in[2][3] = 13;
		pixel_array_in[3][0] = 4;
		pixel_array_in[3][1] = 8;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 33;
		#10;
		
		$display("Input: \n[[35, 26, 43, 9],\n[34, 25, 44, 39],\n[54, 58, 58, 58],\n[21, 5, 53, 17]]");
		$display("Expect: 179, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 43;
		pixel_array_in[0][1] = 42;
		pixel_array_in[0][2] = 54;
		pixel_array_in[0][3] = 55;
		pixel_array_in[1][0] = 41;
		pixel_array_in[1][1] = 17;
		pixel_array_in[1][2] = 9;
		pixel_array_in[1][3] = 16;
		pixel_array_in[2][0] = 44;
		pixel_array_in[2][1] = 29;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 54;
		pixel_array_in[3][1] = 19;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 59;
		#10;
		
		$display("Input: \n[[5, 28, 53, 62],\n[4, 50, 28, 31],\n[33, 32, 33, 60],\n[21, 23, 61, 37]]");
		$display("Expect: 171, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 60;
		pixel_array_in[0][1] = 27;
		pixel_array_in[0][2] = 61;
		pixel_array_in[0][3] = 28;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 21;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 45;
		pixel_array_in[2][0] = 7;
		pixel_array_in[2][1] = 41;
		pixel_array_in[2][2] = 42;
		pixel_array_in[2][3] = 6;
		pixel_array_in[3][0] = 34;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 9;
		pixel_array_in[3][3] = 51;
		#10;
		
		$display("Input: \n[[25, 55, 44, 62],\n[31, 60, 37, 19],\n[6, 53, 6, 13],\n[4, 8, 51, 33]]");
		$display("Expect: 238, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 12;
		pixel_array_in[0][1] = 34;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 46;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 51;
		pixel_array_in[1][2] = 17;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 37;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 29;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 40;
		pixel_array_in[3][2] = 41;
		pixel_array_in[3][3] = 45;
		#10;
		
		$display("Input: \n[[43, 42, 54, 55],\n[41, 17, 9, 16],\n[44, 29, 57, 24],\n[54, 19, 36, 59]]");
		$display("Expect: 88, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 46;
		pixel_array_in[0][1] = 29;
		pixel_array_in[0][2] = 56;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 42;
		pixel_array_in[1][2] = 19;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 19;
		pixel_array_in[2][1] = 21;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 13;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 16;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[60, 27, 61, 28],\n[58, 21, 3, 45],\n[7, 41, 42, 6],\n[34, 18, 9, 51]]");
		$display("Expect: 128, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 18;
		pixel_array_in[0][1] = 33;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 20;
		pixel_array_in[1][0] = 16;
		pixel_array_in[1][1] = 11;
		pixel_array_in[1][2] = 49;
		pixel_array_in[1][3] = 22;
		pixel_array_in[2][0] = 27;
		pixel_array_in[2][1] = 54;
		pixel_array_in[2][2] = 41;
		pixel_array_in[2][3] = 51;
		pixel_array_in[3][0] = 5;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 5;
		pixel_array_in[3][3] = 29;
		#10;
		
		$display("Input: \n[[12, 34, 4, 46],\n[0, 51, 17, 38],\n[37, 32, 29, 39],\n[36, 40, 41, 45]]");
		$display("Expect: 168, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 1;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 27;
		pixel_array_in[1][0] = 7;
		pixel_array_in[1][1] = 58;
		pixel_array_in[1][2] = 36;
		pixel_array_in[1][3] = 45;
		pixel_array_in[2][0] = 12;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 15;
		pixel_array_in[3][0] = 0;
		pixel_array_in[3][1] = 9;
		pixel_array_in[3][2] = 18;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[46, 29, 56, 41],\n[44, 42, 19, 18],\n[19, 21, 19, 13],\n[32, 28, 16, 2]]");
		$display("Expect: 127, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 2;
		pixel_array_in[0][1] = 13;
		pixel_array_in[0][2] = 56;
		pixel_array_in[0][3] = 9;
		pixel_array_in[1][0] = 47;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 56;
		pixel_array_in[1][3] = 55;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 46;
		pixel_array_in[2][2] = 47;
		pixel_array_in[2][3] = 56;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 42;
		pixel_array_in[3][2] = 20;
		pixel_array_in[3][3] = 30;
		#10;
		
		$display("Input: \n[[18, 33, 12, 20],\n[16, 11, 49, 22],\n[27, 54, 41, 51],\n[5, 28, 5, 29]]");
		$display("Expect: 131, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 23;
		pixel_array_in[0][1] = 11;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 35;
		pixel_array_in[1][0] = 11;
		pixel_array_in[1][1] = 61;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 45;
		pixel_array_in[2][0] = 44;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 44;
		pixel_array_in[2][3] = 12;
		pixel_array_in[3][0] = 4;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 17;
		pixel_array_in[3][3] = 28;
		#10;
		
		$display("Input: \n[[53, 1, 30, 27],\n[7, 58, 36, 45],\n[12, 3, 44, 15],\n[0, 9, 18, 6]]");
		$display("Expect: 134, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 15;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 40;
		pixel_array_in[0][3] = 51;
		pixel_array_in[1][0] = 26;
		pixel_array_in[1][1] = 40;
		pixel_array_in[1][2] = 42;
		pixel_array_in[1][3] = 13;
		pixel_array_in[2][0] = 37;
		pixel_array_in[2][1] = 35;
		pixel_array_in[2][2] = 38;
		pixel_array_in[2][3] = 5;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 28;
		pixel_array_in[3][2] = 58;
		pixel_array_in[3][3] = 2;
		#10;
		
		$display("Input: \n[[2, 13, 56, 9],\n[47, 25, 56, 55],\n[30, 46, 47, 56],\n[10, 42, 20, 30]]");
		$display("Expect: 146, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 2;
		pixel_array_in[0][1] = 6;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 52;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 34;
		pixel_array_in[1][2] = 12;
		pixel_array_in[1][3] = 45;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 51;
		pixel_array_in[2][3] = 5;
		pixel_array_in[3][0] = 62;
		pixel_array_in[3][1] = 23;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 5;
		#10;
		
		$display("Input: \n[[23, 11, 32, 35],\n[11, 61, 13, 45],\n[44, 17, 44, 12],\n[4, 25, 17, 28]]");
		$display("Expect: 166, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 2;
		pixel_array_in[0][1] = 38;
		pixel_array_in[0][2] = 61;
		pixel_array_in[0][3] = 6;
		pixel_array_in[1][0] = 50;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 27;
		pixel_array_in[1][3] = 48;
		pixel_array_in[2][0] = 46;
		pixel_array_in[2][1] = 22;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 53;
		pixel_array_in[3][0] = 18;
		pixel_array_in[3][1] = 51;
		pixel_array_in[3][2] = 13;
		pixel_array_in[3][3] = 3;
		#10;
		
		$display("Input: \n[[15, 52, 40, 51],\n[26, 40, 42, 13],\n[37, 35, 38, 5],\n[10, 28, 58, 2]]");
		$display("Expect: 148, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 40;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 58;
		pixel_array_in[0][3] = 38;
		pixel_array_in[1][0] = 39;
		pixel_array_in[1][1] = 31;
		pixel_array_in[1][2] = 48;
		pixel_array_in[1][3] = 43;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 61;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 30;
		pixel_array_in[3][2] = 32;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[2, 6, 48, 52],\n[38, 34, 12, 45],\n[43, 23, 51, 5],\n[62, 23, 11, 5]]");
		$display("Expect: 121, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 49;
		pixel_array_in[0][2] = 39;
		pixel_array_in[0][3] = 58;
		pixel_array_in[1][0] = 62;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 16;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 56;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 34;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[2, 38, 61, 6],\n[50, 7, 27, 48],\n[46, 22, 7, 53],\n[18, 51, 13, 3]]");
		$display("Expect: 43, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 17;
		pixel_array_in[0][1] = 19;
		pixel_array_in[0][2] = 43;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 61;
		pixel_array_in[1][1] = 31;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 54;
		pixel_array_in[2][0] = 61;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 41;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 62;
		pixel_array_in[3][3] = 48;
		#10;
		
		$display("Input: \n[[40, 56, 58, 38],\n[39, 31, 48, 43],\n[22, 61, 23, 9],\n[32, 30, 32, 56]]");
		$display("Expect: 185, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 46;
		pixel_array_in[0][1] = 34;
		pixel_array_in[0][2] = 1;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 9;
		pixel_array_in[1][2] = 45;
		pixel_array_in[1][3] = 36;
		pixel_array_in[2][0] = 22;
		pixel_array_in[2][1] = 21;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 31;
		pixel_array_in[3][0] = 50;
		pixel_array_in[3][1] = 47;
		pixel_array_in[3][2] = 51;
		pixel_array_in[3][3] = 54;
		#10;
		
		$display("Input: \n[[0, 49, 39, 58],\n[62, 7, 16, 46],\n[15, 56, 49, 55],\n[34, 34, 29, 35]]");
		$display("Expect: 121, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 21;
		pixel_array_in[0][1] = 32;
		pixel_array_in[0][2] = 59;
		pixel_array_in[0][3] = 11;
		pixel_array_in[1][0] = 13;
		pixel_array_in[1][1] = 54;
		pixel_array_in[1][2] = 32;
		pixel_array_in[1][3] = 54;
		pixel_array_in[2][0] = 52;
		pixel_array_in[2][1] = 20;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 56;
		pixel_array_in[3][1] = 22;
		pixel_array_in[3][2] = 10;
		pixel_array_in[3][3] = 6;
		#10;
		
		$display("Input: \n[[17, 19, 43, 42],\n[61, 31, 22, 54],\n[61, 17, 41, 25],\n[42, 25, 62, 48]]");
		$display("Expect: 97, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 33;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 51;
		pixel_array_in[1][0] = 3;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 3;
		pixel_array_in[1][3] = 36;
		pixel_array_in[2][0] = 30;
		pixel_array_in[2][1] = 46;
		pixel_array_in[2][2] = 27;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 11;
		pixel_array_in[3][1] = 62;
		pixel_array_in[3][2] = 38;
		pixel_array_in[3][3] = 3;
		#10;
		
		$display("Input: \n[[46, 34, 1, 42],\n[58, 9, 45, 36],\n[22, 21, 49, 31],\n[50, 47, 51, 54]]");
		$display("Expect: 47, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 6;
		pixel_array_in[0][1] = 25;
		pixel_array_in[0][2] = 9;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 0;
		pixel_array_in[1][1] = 26;
		pixel_array_in[1][2] = 59;
		pixel_array_in[1][3] = 13;
		pixel_array_in[2][0] = 40;
		pixel_array_in[2][1] = 61;
		pixel_array_in[2][2] = 36;
		pixel_array_in[2][3] = 52;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 50;
		pixel_array_in[3][3] = 22;
		#10;
		
		$display("Input: \n[[21, 32, 59, 11],\n[13, 54, 32, 54],\n[52, 20, 19, 43],\n[56, 22, 10, 6]]");
		$display("Expect: 153, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 8;
		pixel_array_in[0][1] = 61;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 23;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 37;
		pixel_array_in[1][2] = 57;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 48;
		pixel_array_in[2][2] = 19;
		pixel_array_in[2][3] = 33;
		pixel_array_in[3][0] = 42;
		pixel_array_in[3][1] = 2;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[33, 7, 48, 51],\n[3, 50, 3, 36],\n[30, 46, 27, 24],\n[11, 62, 38, 3]]");
		$display("Expect: 198, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 4;
		pixel_array_in[0][2] = 15;
		pixel_array_in[0][3] = 50;
		pixel_array_in[1][0] = 46;
		pixel_array_in[1][1] = 42;
		pixel_array_in[1][2] = 16;
		pixel_array_in[1][3] = 30;
		pixel_array_in[2][0] = 13;
		pixel_array_in[2][1] = 32;
		pixel_array_in[2][2] = 52;
		pixel_array_in[2][3] = 33;
		pixel_array_in[3][0] = 16;
		pixel_array_in[3][1] = 5;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 50;
		#10;
		
		$display("Input: \n[[6, 25, 9, 57],\n[0, 26, 59, 13],\n[40, 61, 36, 52],\n[32, 34, 50, 22]]");
		$display("Expect: 181, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 22;
		pixel_array_in[0][1] = 51;
		pixel_array_in[0][2] = 61;
		pixel_array_in[0][3] = 33;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 57;
		pixel_array_in[1][2] = 52;
		pixel_array_in[1][3] = 51;
		pixel_array_in[2][0] = 3;
		pixel_array_in[2][1] = 25;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 59;
		pixel_array_in[3][1] = 52;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 30;
		#10;
		
		$display("Input: \n[[8, 61, 34, 23],\n[22, 37, 57, 0],\n[57, 48, 19, 33],\n[42, 2, 11, 35]]");
		$display("Expect: 175, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 59;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 5;
		pixel_array_in[0][3] = 46;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 61;
		pixel_array_in[1][2] = 7;
		pixel_array_in[1][3] = 59;
		pixel_array_in[2][0] = 62;
		pixel_array_in[2][1] = 44;
		pixel_array_in[2][2] = 1;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 37;
		pixel_array_in[3][1] = 56;
		pixel_array_in[3][2] = 20;
		pixel_array_in[3][3] = 61;
		#10;
		
		$display("Input: \n[[19, 4, 15, 50],\n[46, 42, 16, 30],\n[13, 32, 52, 33],\n[16, 5, 27, 50]]");
		$display("Expect: 164, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 23;
		pixel_array_in[0][2] = 7;
		pixel_array_in[0][3] = 49;
		pixel_array_in[1][0] = 1;
		pixel_array_in[1][1] = 50;
		pixel_array_in[1][2] = 22;
		pixel_array_in[1][3] = 27;
		pixel_array_in[2][0] = 37;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 31;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 61;
		pixel_array_in[3][3] = 50;
		#10;
		
		$display("Input: \n[[22, 51, 61, 33],\n[31, 57, 52, 51],\n[3, 25, 54, 9],\n[59, 52, 29, 30]]");
		$display("Expect: 158, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 35;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 54;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 9;
		pixel_array_in[1][1] = 52;
		pixel_array_in[1][2] = 7;
		pixel_array_in[1][3] = 49;
		pixel_array_in[2][0] = 59;
		pixel_array_in[2][1] = 29;
		pixel_array_in[2][2] = 48;
		pixel_array_in[2][3] = 22;
		pixel_array_in[3][0] = 52;
		pixel_array_in[3][1] = 45;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[59, 18, 5, 46],\n[32, 61, 7, 59],\n[62, 44, 1, 44],\n[37, 56, 20, 61]]");
		$display("Expect: 217, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 58;
		pixel_array_in[0][1] = 56;
		pixel_array_in[0][2] = 10;
		pixel_array_in[0][3] = 14;
		pixel_array_in[1][0] = 38;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 35;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 53;
		pixel_array_in[2][2] = 3;
		pixel_array_in[2][3] = 29;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[19, 23, 7, 49],\n[1, 50, 22, 27],\n[37, 17, 31, 24],\n[52, 48, 61, 50]]");
		$display("Expect: 133, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 7;
		pixel_array_in[0][1] = 15;
		pixel_array_in[0][2] = 42;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 30;
		pixel_array_in[1][1] = 48;
		pixel_array_in[1][2] = 42;
		pixel_array_in[1][3] = 47;
		pixel_array_in[2][0] = 20;
		pixel_array_in[2][1] = 58;
		pixel_array_in[2][2] = 10;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 6;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 15;
		pixel_array_in[3][3] = 9;
		#10;
		
		$display("Input: \n[[35, 7, 54, 2],\n[9, 52, 7, 49],\n[59, 29, 48, 22],\n[52, 45, 48, 35]]");
		$display("Expect: 169, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 0;
		pixel_array_in[0][1] = 53;
		pixel_array_in[0][2] = 18;
		pixel_array_in[0][3] = 37;
		pixel_array_in[1][0] = 12;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 6;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 46;
		pixel_array_in[2][1] = 4;
		pixel_array_in[2][2] = 0;
		pixel_array_in[2][3] = 35;
		pixel_array_in[3][0] = 48;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 9;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[58, 56, 10, 14],\n[38, 35, 35, 15],\n[50, 53, 3, 29],\n[25, 6, 60, 1]]");
		$display("Expect: 182, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 40;
		pixel_array_in[0][1] = 38;
		pixel_array_in[0][2] = 48;
		pixel_array_in[0][3] = 45;
		pixel_array_in[1][0] = 32;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 25;
		pixel_array_in[1][3] = 43;
		pixel_array_in[2][0] = 52;
		pixel_array_in[2][1] = 37;
		pixel_array_in[2][2] = 59;
		pixel_array_in[2][3] = 8;
		pixel_array_in[3][0] = 51;
		pixel_array_in[3][1] = 0;
		pixel_array_in[3][2] = 39;
		pixel_array_in[3][3] = 7;
		#10;
		
		$display("Input: \n[[7, 15, 42, 25],\n[30, 48, 42, 47],\n[20, 58, 10, 32],\n[6, 58, 15, 9]]");
		$display("Expect: 220, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 48;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 53;
		pixel_array_in[0][3] = 41;
		pixel_array_in[1][0] = 53;
		pixel_array_in[1][1] = 60;
		pixel_array_in[1][2] = 18;
		pixel_array_in[1][3] = 32;
		pixel_array_in[2][0] = 53;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 52;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 14;
		pixel_array_in[3][2] = 35;
		pixel_array_in[3][3] = 19;
		#10;
		
		$display("Input: \n[[0, 53, 18, 37],\n[12, 27, 6, 35],\n[46, 4, 0, 35],\n[48, 0, 9, 52]]");
		$display("Expect: 56, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 9;
		pixel_array_in[0][1] = 12;
		pixel_array_in[0][2] = 34;
		pixel_array_in[0][3] = 34;
		pixel_array_in[1][0] = 25;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 34;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 42;
		pixel_array_in[2][1] = 8;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 28;
		pixel_array_in[3][1] = 8;
		pixel_array_in[3][2] = 27;
		pixel_array_in[3][3] = 30;
		#10;
		
		$display("Input: \n[[40, 38, 48, 45],\n[32, 12, 25, 43],\n[52, 37, 59, 8],\n[51, 0, 39, 7]]");
		$display("Expect: 100, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 13;
		pixel_array_in[0][1] = 21;
		pixel_array_in[0][2] = 30;
		pixel_array_in[0][3] = 38;
		pixel_array_in[1][0] = 1;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 27;
		pixel_array_in[1][3] = 44;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 23;
		pixel_array_in[2][2] = 29;
		pixel_array_in[2][3] = 2;
		pixel_array_in[3][0] = 27;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 21;
		#10;
		
		$display("Input: \n[[48, 18, 53, 41],\n[53, 60, 18, 32],\n[53, 3, 61, 52],\n[10, 14, 35, 19]]");
		$display("Expect: 133, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 18;
		pixel_array_in[0][1] = 9;
		pixel_array_in[0][2] = 50;
		pixel_array_in[0][3] = 8;
		pixel_array_in[1][0] = 42;
		pixel_array_in[1][1] = 33;
		pixel_array_in[1][2] = 40;
		pixel_array_in[1][3] = 17;
		pixel_array_in[2][0] = 43;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 22;
		pixel_array_in[2][3] = 39;
		pixel_array_in[3][0] = 37;
		pixel_array_in[3][1] = 50;
		pixel_array_in[3][2] = 57;
		pixel_array_in[3][3] = 42;
		#10;
		
		$display("Input: \n[[9, 12, 34, 34],\n[25, 23, 34, 38],\n[42, 8, 23, 3],\n[28, 8, 27, 30]]");
		$display("Expect: 64, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 47;
		pixel_array_in[0][1] = 5;
		pixel_array_in[0][2] = 2;
		pixel_array_in[0][3] = 49;
		pixel_array_in[1][0] = 4;
		pixel_array_in[1][1] = 19;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 49;
		pixel_array_in[2][0] = 34;
		pixel_array_in[2][1] = 46;
		pixel_array_in[2][2] = 7;
		pixel_array_in[2][3] = 9;
		pixel_array_in[3][0] = 59;
		pixel_array_in[3][1] = 21;
		pixel_array_in[3][2] = 8;
		pixel_array_in[3][3] = 56;
		#10;
		
		$display("Input: \n[[13, 21, 30, 38],\n[1, 7, 27, 44],\n[57, 23, 29, 2],\n[27, 34, 7, 21]]");
		$display("Expect: 53, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 24;
		pixel_array_in[0][1] = 28;
		pixel_array_in[0][2] = 3;
		pixel_array_in[0][3] = 50;
		pixel_array_in[1][0] = 2;
		pixel_array_in[1][1] = 18;
		pixel_array_in[1][2] = 1;
		pixel_array_in[1][3] = 1;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 37;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 34;
		pixel_array_in[3][2] = 43;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[18, 9, 50, 8],\n[42, 33, 40, 17],\n[43, 17, 22, 39],\n[37, 50, 57, 42]]");
		$display("Expect: 97, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 39;
		pixel_array_in[0][1] = 30;
		pixel_array_in[0][2] = 13;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 44;
		pixel_array_in[1][1] = 26;
		pixel_array_in[1][2] = 38;
		pixel_array_in[1][3] = 9;
		pixel_array_in[2][0] = 56;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 33;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 61;
		pixel_array_in[3][1] = 58;
		pixel_array_in[3][2] = 2;
		pixel_array_in[3][3] = 27;
		#10;
		
		$display("Input: \n[[47, 5, 2, 49],\n[4, 19, 13, 49],\n[34, 46, 7, 9],\n[59, 21, 8, 56]]");
		$display("Expect: 139, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 6;
		pixel_array_in[0][1] = 57;
		pixel_array_in[0][2] = 39;
		pixel_array_in[0][3] = 15;
		pixel_array_in[1][0] = 42;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 54;
		pixel_array_in[1][3] = 1;
		pixel_array_in[2][0] = 58;
		pixel_array_in[2][1] = 49;
		pixel_array_in[2][2] = 26;
		pixel_array_in[2][3] = 56;
		pixel_array_in[3][0] = 43;
		pixel_array_in[3][1] = 33;
		pixel_array_in[3][2] = 7;
		pixel_array_in[3][3] = 44;
		#10;
		
		$display("Input: \n[[24, 28, 3, 50],\n[2, 18, 1, 1],\n[1, 13, 37, 44],\n[19, 34, 43, 39]]");
		$display("Expect: 54, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 39;
		pixel_array_in[0][1] = 54;
		pixel_array_in[0][2] = 25;
		pixel_array_in[0][3] = 40;
		pixel_array_in[1][0] = 28;
		pixel_array_in[1][1] = 3;
		pixel_array_in[1][2] = 14;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 28;
		pixel_array_in[2][1] = 25;
		pixel_array_in[2][2] = 39;
		pixel_array_in[2][3] = 60;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 47;
		pixel_array_in[3][2] = 45;
		pixel_array_in[3][3] = 28;
		#10;
		
		$display("Input: \n[[39, 30, 13, 59],\n[44, 26, 38, 9],\n[56, 7, 33, 55],\n[61, 58, 2, 27]]");
		$display("Expect: 52, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 14;
		pixel_array_in[0][1] = 42;
		pixel_array_in[0][2] = 19;
		pixel_array_in[0][3] = 54;
		pixel_array_in[1][0] = 48;
		pixel_array_in[1][1] = 56;
		pixel_array_in[1][2] = 29;
		pixel_array_in[1][3] = 36;
		pixel_array_in[2][0] = 59;
		pixel_array_in[2][1] = 22;
		pixel_array_in[2][2] = 48;
		pixel_array_in[2][3] = 18;
		pixel_array_in[3][0] = 32;
		pixel_array_in[3][1] = 51;
		pixel_array_in[3][2] = 4;
		pixel_array_in[3][3] = 46;
		#10;
		
		$display("Input: \n[[6, 57, 39, 15],\n[42, 25, 54, 1],\n[58, 49, 26, 56],\n[43, 33, 7, 44]]");
		$display("Expect: 144, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 26;
		pixel_array_in[0][1] = 51;
		pixel_array_in[0][2] = 8;
		pixel_array_in[0][3] = 51;
		pixel_array_in[1][0] = 33;
		pixel_array_in[1][1] = 25;
		pixel_array_in[1][2] = 50;
		pixel_array_in[1][3] = 15;
		pixel_array_in[2][0] = 10;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 57;
		pixel_array_in[2][3] = 24;
		pixel_array_in[3][0] = 33;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 31;
		pixel_array_in[3][3] = 8;
		#10;
		
		$display("Input: \n[[39, 54, 25, 40],\n[28, 3, 14, 15],\n[28, 25, 39, 60],\n[19, 47, 45, 28]]");
		$display("Expect: 37, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 53;
		pixel_array_in[0][1] = 52;
		pixel_array_in[0][2] = 4;
		pixel_array_in[0][3] = 3;
		pixel_array_in[1][0] = 33;
		pixel_array_in[1][1] = 23;
		pixel_array_in[1][2] = 34;
		pixel_array_in[1][3] = 18;
		pixel_array_in[2][0] = 61;
		pixel_array_in[2][1] = 19;
		pixel_array_in[2][2] = 43;
		pixel_array_in[2][3] = 45;
		pixel_array_in[3][0] = 13;
		pixel_array_in[3][1] = 47;
		pixel_array_in[3][2] = 44;
		pixel_array_in[3][3] = 1;
		#10;
		
		$display("Input: \n[[14, 42, 19, 54],\n[48, 56, 29, 36],\n[59, 22, 48, 18],\n[32, 51, 4, 46]]");
		$display("Expect: 152, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 19;
		pixel_array_in[0][1] = 43;
		pixel_array_in[0][2] = 27;
		pixel_array_in[0][3] = 1;
		pixel_array_in[1][0] = 24;
		pixel_array_in[1][1] = 22;
		pixel_array_in[1][2] = 41;
		pixel_array_in[1][3] = 55;
		pixel_array_in[2][0] = 59;
		pixel_array_in[2][1] = 22;
		pixel_array_in[2][2] = 32;
		pixel_array_in[2][3] = 44;
		pixel_array_in[3][0] = 25;
		pixel_array_in[3][1] = 25;
		pixel_array_in[3][2] = 49;
		pixel_array_in[3][3] = 46;
		#10;
		
		$display("Input: \n[[26, 51, 8, 51],\n[33, 25, 50, 15],\n[10, 17, 57, 24],\n[33, 6, 31, 8]]");
		$display("Expect: 80, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 59;
		pixel_array_in[0][1] = 2;
		pixel_array_in[0][2] = 6;
		pixel_array_in[0][3] = 57;
		pixel_array_in[1][0] = 19;
		pixel_array_in[1][1] = 57;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 35;
		pixel_array_in[2][0] = 55;
		pixel_array_in[2][1] = 39;
		pixel_array_in[2][2] = 61;
		pixel_array_in[2][3] = 32;
		pixel_array_in[3][0] = 24;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 57;
		pixel_array_in[3][3] = 52;
		#10;
		
		$display("Input: \n[[53, 52, 4, 3],\n[33, 23, 34, 18],\n[61, 19, 43, 45],\n[13, 47, 44, 1]]");
		$display("Expect: 69, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 44;
		pixel_array_in[0][1] = 15;
		pixel_array_in[0][2] = 32;
		pixel_array_in[0][3] = 56;
		pixel_array_in[1][0] = 41;
		pixel_array_in[1][1] = 49;
		pixel_array_in[1][2] = 33;
		pixel_array_in[1][3] = 4;
		pixel_array_in[2][0] = 26;
		pixel_array_in[2][1] = 10;
		pixel_array_in[2][2] = 24;
		pixel_array_in[2][3] = 50;
		pixel_array_in[3][0] = 11;
		pixel_array_in[3][1] = 12;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 39;
		#10;
		
		$display("Input: \n[[19, 43, 27, 1],\n[24, 22, 41, 55],\n[59, 22, 32, 44],\n[25, 25, 49, 46]]");
		$display("Expect: 82, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 1;
		pixel_array_in[0][1] = 34;
		pixel_array_in[0][2] = 12;
		pixel_array_in[0][3] = 51;
		pixel_array_in[1][0] = 18;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 18;
		pixel_array_in[1][3] = 41;
		pixel_array_in[2][0] = 52;
		pixel_array_in[2][1] = 3;
		pixel_array_in[2][2] = 15;
		pixel_array_in[2][3] = 46;
		pixel_array_in[3][0] = 31;
		pixel_array_in[3][1] = 6;
		pixel_array_in[3][2] = 59;
		pixel_array_in[3][3] = 4;
		#10;
		
		$display("Input: \n[[59, 2, 6, 57],\n[19, 57, 33, 35],\n[55, 39, 61, 32],\n[24, 37, 57, 52]]");
		$display("Expect: 206, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 41;
		pixel_array_in[0][1] = 48;
		pixel_array_in[0][2] = 37;
		pixel_array_in[0][3] = 25;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 12;
		pixel_array_in[1][2] = 59;
		pixel_array_in[1][3] = 13;
		pixel_array_in[2][0] = 50;
		pixel_array_in[2][1] = 14;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 3;
		pixel_array_in[3][0] = 36;
		pixel_array_in[3][1] = 18;
		pixel_array_in[3][2] = 6;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[44, 15, 32, 56],\n[41, 49, 33, 4],\n[26, 10, 24, 50],\n[11, 12, 48, 39]]");
		$display("Expect: 126, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 35;
		pixel_array_in[0][1] = 49;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 42;
		pixel_array_in[1][0] = 49;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 49;
		pixel_array_in[1][3] = 53;
		pixel_array_in[2][0] = 9;
		pixel_array_in[2][1] = 2;
		pixel_array_in[2][2] = 31;
		pixel_array_in[2][3] = 14;
		pixel_array_in[3][0] = 55;
		pixel_array_in[3][1] = 43;
		pixel_array_in[3][2] = 11;
		pixel_array_in[3][3] = 41;
		#10;
		
		$display("Input: \n[[1, 34, 12, 51],\n[18, 12, 18, 41],\n[52, 3, 15, 46],\n[31, 6, 59, 4]]");
		$display("Expect: 23, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 7;
		pixel_array_in[0][2] = 28;
		pixel_array_in[0][3] = 22;
		pixel_array_in[1][0] = 17;
		pixel_array_in[1][1] = 27;
		pixel_array_in[1][2] = 17;
		pixel_array_in[1][3] = 56;
		pixel_array_in[2][0] = 27;
		pixel_array_in[2][1] = 17;
		pixel_array_in[2][2] = 26;
		pixel_array_in[2][3] = 26;
		pixel_array_in[3][0] = 2;
		pixel_array_in[3][1] = 52;
		pixel_array_in[3][2] = 29;
		pixel_array_in[3][3] = 16;
		#10;
		
		$display("Input: \n[[41, 48, 37, 25],\n[58, 12, 59, 13],\n[50, 14, 5, 3],\n[36, 18, 6, 16]]");
		$display("Expect: 42, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 54;
		pixel_array_in[0][1] = 15;
		pixel_array_in[0][2] = 55;
		pixel_array_in[0][3] = 2;
		pixel_array_in[1][0] = 34;
		pixel_array_in[1][1] = 22;
		pixel_array_in[1][2] = 53;
		pixel_array_in[1][3] = 46;
		pixel_array_in[2][0] = 51;
		pixel_array_in[2][1] = 12;
		pixel_array_in[2][2] = 23;
		pixel_array_in[2][3] = 31;
		pixel_array_in[3][0] = 28;
		pixel_array_in[3][1] = 56;
		pixel_array_in[3][2] = 16;
		pixel_array_in[3][3] = 5;
		#10;
		
		$display("Input: \n[[35, 49, 45, 42],\n[49, 45, 49, 53],\n[9, 2, 31, 14],\n[55, 43, 11, 41]]");
		$display("Expect: 82, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 60;
		pixel_array_in[0][1] = 61;
		pixel_array_in[0][2] = 56;
		pixel_array_in[0][3] = 27;
		pixel_array_in[1][0] = 58;
		pixel_array_in[1][1] = 32;
		pixel_array_in[1][2] = 35;
		pixel_array_in[1][3] = 53;
		pixel_array_in[2][0] = 9;
		pixel_array_in[2][1] = 37;
		pixel_array_in[2][2] = 49;
		pixel_array_in[2][3] = 25;
		pixel_array_in[3][0] = 11;
		pixel_array_in[3][1] = 38;
		pixel_array_in[3][2] = 53;
		pixel_array_in[3][3] = 3;
		#10;
		
		$display("Input: \n[[61, 7, 28, 22],\n[17, 27, 17, 56],\n[27, 17, 26, 26],\n[2, 52, 29, 16]]");
		$display("Expect: 84, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 35;
		pixel_array_in[0][1] = 15;
		pixel_array_in[0][2] = 23;
		pixel_array_in[0][3] = 30;
		pixel_array_in[1][0] = 31;
		pixel_array_in[1][1] = 21;
		pixel_array_in[1][2] = 39;
		pixel_array_in[1][3] = 5;
		pixel_array_in[2][0] = 58;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 24;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 19;
		pixel_array_in[3][1] = 15;
		pixel_array_in[3][2] = 28;
		pixel_array_in[3][3] = 58;
		#10;
		
		$display("Input: \n[[54, 15, 55, 2],\n[34, 22, 53, 46],\n[51, 12, 23, 31],\n[28, 56, 16, 5]]");
		$display("Expect: 58, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 43;
		pixel_array_in[0][1] = 46;
		pixel_array_in[0][2] = 8;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 24;
		pixel_array_in[1][1] = 26;
		pixel_array_in[1][2] = 26;
		pixel_array_in[1][3] = 33;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 42;
		pixel_array_in[2][2] = 16;
		pixel_array_in[2][3] = 43;
		pixel_array_in[3][0] = 29;
		pixel_array_in[3][1] = 9;
		pixel_array_in[3][2] = 4;
		pixel_array_in[3][3] = 18;
		#10;
		
		$display("Input: \n[[60, 61, 56, 27],\n[58, 32, 35, 53],\n[9, 37, 49, 25],\n[11, 38, 53, 3]]");
		$display("Expect: 130, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 34;
		pixel_array_in[0][1] = 16;
		pixel_array_in[0][2] = 6;
		pixel_array_in[0][3] = 47;
		pixel_array_in[1][0] = 16;
		pixel_array_in[1][1] = 7;
		pixel_array_in[1][2] = 44;
		pixel_array_in[1][3] = 38;
		pixel_array_in[2][0] = 14;
		pixel_array_in[2][1] = 56;
		pixel_array_in[2][2] = 45;
		pixel_array_in[2][3] = 30;
		pixel_array_in[3][0] = 6;
		pixel_array_in[3][1] = 1;
		pixel_array_in[3][2] = 48;
		pixel_array_in[3][3] = 62;
		#10;
		
		$display("Input: \n[[35, 15, 23, 30],\n[31, 21, 39, 5],\n[58, 7, 24, 30],\n[19, 15, 28, 58]]");
		$display("Expect: 55, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 49;
		pixel_array_in[0][1] = 38;
		pixel_array_in[0][2] = 9;
		pixel_array_in[0][3] = 13;
		pixel_array_in[1][0] = 22;
		pixel_array_in[1][1] = 35;
		pixel_array_in[1][2] = 12;
		pixel_array_in[1][3] = 21;
		pixel_array_in[2][0] = 15;
		pixel_array_in[2][1] = 59;
		pixel_array_in[2][2] = 55;
		pixel_array_in[2][3] = 49;
		pixel_array_in[3][0] = 15;
		pixel_array_in[3][1] = 48;
		pixel_array_in[3][2] = 34;
		pixel_array_in[3][3] = 35;
		#10;
		
		$display("Input: \n[[43, 46, 8, 59],\n[24, 26, 26, 33],\n[1, 42, 16, 43],\n[29, 9, 4, 18]]");
		$display("Expect: 139, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 61;
		pixel_array_in[0][1] = 43;
		pixel_array_in[0][2] = 50;
		pixel_array_in[0][3] = 59;
		pixel_array_in[1][0] = 23;
		pixel_array_in[1][1] = 43;
		pixel_array_in[1][2] = 61;
		pixel_array_in[1][3] = 3;
		pixel_array_in[2][0] = 1;
		pixel_array_in[2][1] = 53;
		pixel_array_in[2][2] = 54;
		pixel_array_in[2][3] = 52;
		pixel_array_in[3][0] = 46;
		pixel_array_in[3][1] = 37;
		pixel_array_in[3][2] = 60;
		pixel_array_in[3][3] = 32;
		#10;
		
		$display("Input: \n[[34, 16, 6, 47],\n[16, 7, 44, 38],\n[14, 56, 45, 30],\n[6, 1, 48, 62]]");
		$display("Expect: 137, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 33;
		pixel_array_in[0][1] = 22;
		pixel_array_in[0][2] = 2;
		pixel_array_in[0][3] = 46;
		pixel_array_in[1][0] = 55;
		pixel_array_in[1][1] = 2;
		pixel_array_in[1][2] = 13;
		pixel_array_in[1][3] = 49;
		pixel_array_in[2][0] = 57;
		pixel_array_in[2][1] = 13;
		pixel_array_in[2][2] = 5;
		pixel_array_in[2][3] = 55;
		pixel_array_in[3][0] = 10;
		pixel_array_in[3][1] = 32;
		pixel_array_in[3][2] = 8;
		pixel_array_in[3][3] = 50;
		#10;
		
		$display("Input: \n[[49, 38, 9, 13],\n[22, 35, 12, 21],\n[15, 59, 55, 49],\n[15, 48, 34, 35]]");
		$display("Expect: 190, Result: %d", pixel_out);
		$display("");
		pixel_array_in[0][0] = 18;
		pixel_array_in[0][1] = 18;
		pixel_array_in[0][2] = 45;
		pixel_array_in[0][3] = 26;
		pixel_array_in[1][0] = 18;
		pixel_array_in[1][1] = 45;
		pixel_array_in[1][2] = 45;
		pixel_array_in[1][3] = 0;
		pixel_array_in[2][0] = 59;
		pixel_array_in[2][1] = 7;
		pixel_array_in[2][2] = 13;
		pixel_array_in[2][3] = 20;
		pixel_array_in[3][0] = 50;
		pixel_array_in[3][1] = 13;
		pixel_array_in[3][2] = 36;
		pixel_array_in[3][3] = 10;
		#10;
		
		$display("Input: \n[[61, 43, 50, 59],\n[23, 43, 61, 3],\n[1, 53, 54, 52],\n[46, 37, 60, 32]]");
		$display("Expect: 196, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[33, 22, 2, 46],\n[55, 2, 13, 49],\n[57, 13, 5, 55],\n[10, 32, 8, 50]]");
		$display("Expect: 20, Result: %d", pixel_out);
		$display("");
		#10;
		
		$display("Input: \n[[18, 18, 45, 26],\n[18, 45, 45, 0],\n[59, 7, 13, 20],\n[50, 13, 36, 10]]");
		$display("Expect: 109, Result: %d", pixel_out);
		$display("");
		#10;
		
		
		$display("Finishing Sim"); //print nice message
		$finish;
		
    end
endmodule //counter_tb

`default_nettype wire